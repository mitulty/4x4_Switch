-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_1_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_1_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_1_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_1_Daemon;
architecture inputPort_1_Daemon_arch of inputPort_1_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_1_Daemon_CP_3_start: Boolean;
  signal inputPort_1_Daemon_CP_3_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_72_branch_req_0 : boolean;
  signal phi_stmt_82_req_1 : boolean;
  signal phi_stmt_82_req_0 : boolean;
  signal phi_stmt_74_req_0 : boolean;
  signal phi_stmt_74_req_1 : boolean;
  signal phi_stmt_74_ack_0 : boolean;
  signal next_count_down_111_76_buf_req_0 : boolean;
  signal next_count_down_111_76_buf_ack_0 : boolean;
  signal next_count_down_111_76_buf_req_1 : boolean;
  signal next_count_down_111_76_buf_ack_1 : boolean;
  signal RPIPE_in_data_1_81_inst_req_0 : boolean;
  signal RPIPE_in_data_1_81_inst_ack_0 : boolean;
  signal RPIPE_in_data_1_81_inst_req_1 : boolean;
  signal RPIPE_in_data_1_81_inst_ack_1 : boolean;
  signal phi_stmt_82_ack_0 : boolean;
  signal next_last_dest_id_117_85_buf_req_0 : boolean;
  signal next_last_dest_id_117_85_buf_ack_0 : boolean;
  signal next_last_dest_id_117_85_buf_req_1 : boolean;
  signal next_last_dest_id_117_85_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_1_129_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_129_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_129_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_1_129_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_2_138_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_2_138_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_2_138_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_2_138_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_3_147_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_3_147_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_3_147_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_3_147_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_4_156_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_4_156_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_4_156_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_4_156_inst_ack_1 : boolean;
  signal do_while_stmt_72_branch_ack_0 : boolean;
  signal do_while_stmt_72_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_1_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_1_Daemon_CP_3_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_1_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_1_Daemon_CP_3: Block -- control-path 
    signal inputPort_1_Daemon_CP_3_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_1_Daemon_CP_3_elements(0) <= inputPort_1_Daemon_CP_3_start;
    inputPort_1_Daemon_CP_3_symbol <= inputPort_1_Daemon_CP_3_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_71/$entry
      -- CP-element group 0: 	 branch_block_stmt_71/branch_block_stmt_71__entry__
      -- CP-element group 0: 	 branch_block_stmt_71/do_while_stmt_72__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_71/$exit
      -- CP-element group 1: 	 branch_block_stmt_71/branch_block_stmt_71__exit__
      -- CP-element group 1: 	 branch_block_stmt_71/do_while_stmt_72__exit__
      -- 
    inputPort_1_Daemon_CP_3_elements(1) <= inputPort_1_Daemon_CP_3_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_71/do_while_stmt_72/$entry
      -- CP-element group 2: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72__entry__
      -- 
    inputPort_1_Daemon_CP_3_elements(2) <= inputPort_1_Daemon_CP_3_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72__exit__
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_71/do_while_stmt_72/loop_back
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	70 
    -- CP-element group 5: 	71 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_71/do_while_stmt_72/condition_done
      -- CP-element group 5: 	 branch_block_stmt_71/do_while_stmt_72/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_71/do_while_stmt_72/loop_taken/$entry
      -- 
    inputPort_1_Daemon_CP_3_elements(5) <= inputPort_1_Daemon_CP_3_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_71/do_while_stmt_72/loop_body_done
      -- 
    inputPort_1_Daemon_CP_3_elements(6) <= inputPort_1_Daemon_CP_3_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/back_edge_to_loop_body
      -- 
    inputPort_1_Daemon_CP_3_elements(7) <= inputPort_1_Daemon_CP_3_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/first_time_through_loop_body
      -- 
    inputPort_1_Daemon_CP_3_elements(8) <= inputPort_1_Daemon_CP_3_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	68 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_79_sample_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/condition_evaluated
      -- 
    condition_evaluated_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(10), ack => do_while_stmt_72_branch_req_0); -- 
    inputPort_1_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(14) & inputPort_1_Daemon_CP_3_elements(68);
      gj_inputPort_1_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_sample_start__ps
      -- 
    inputPort_1_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(15) & inputPort_1_Daemon_CP_3_elements(37) & inputPort_1_Daemon_CP_3_elements(14);
      gj_inputPort_1_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_79_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_sample_completed_
      -- 
    inputPort_1_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(17) & inputPort_1_Daemon_CP_3_elements(35) & inputPort_1_Daemon_CP_3_elements(40);
      gj_inputPort_1_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_update_start__ps
      -- 
    inputPort_1_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(16) & inputPort_1_Daemon_CP_3_elements(32) & inputPort_1_Daemon_CP_3_elements(38);
      gj_inputPort_1_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_1_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42);
      gj_inputPort_1_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_sample_start_
      -- 
    inputPort_1_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(12);
      gj_inputPort_1_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(60) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(66);
      gj_inputPort_1_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_loopback_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(19) <= inputPort_1_Daemon_CP_3_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_loopback_sample_req_ps
      -- 
    phi_stmt_74_loopback_sample_req_42_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_74_loopback_sample_req_42_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(20), ack => phi_stmt_74_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_entry_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(21) <= inputPort_1_Daemon_CP_3_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_entry_sample_req_ps
      -- 
    phi_stmt_74_entry_sample_req_45_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_74_entry_sample_req_45_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(22), ack => phi_stmt_74_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_74_phi_mux_ack_ps
      -- 
    phi_stmt_74_phi_mux_ack_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_74_ack_0, ack => inputPort_1_Daemon_CP_3_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_Sample/req
      -- 
    req_61_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_61_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(24), ack => next_count_down_111_76_buf_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_update_start_
      -- CP-element group 25: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_Update/req
      -- 
    req_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(25), ack => next_count_down_111_76_buf_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_Sample/ack
      -- 
    ack_62_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_111_76_buf_ack_0, ack => inputPort_1_Daemon_CP_3_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_count_down_76_Update/ack
      -- 
    ack_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_111_76_buf_ack_1, ack => inputPort_1_Daemon_CP_3_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/type_cast_78_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/type_cast_78_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/type_cast_78_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/type_cast_78_sample_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/type_cast_78_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/type_cast_78_update_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/type_cast_78_update_completed__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(30) <= inputPort_1_Daemon_CP_3_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/type_cast_78_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(29), ack => inputPort_1_Daemon_CP_3_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_79_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(60) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(66);
      gj_inputPort_1_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_Sample/rr
      -- 
    rr_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(33), ack => RPIPE_in_data_1_81_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(11) & inputPort_1_Daemon_CP_3_elements(36);
      gj_inputPort_1_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_update_start_
      -- CP-element group 34: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_Update/cr
      -- 
    cr_93_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_93_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(34), ack => RPIPE_in_data_1_81_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(13) & inputPort_1_Daemon_CP_3_elements(35);
      gj_inputPort_1_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_Sample/ra
      -- 
    ra_89_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1_81_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_79_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/RPIPE_in_data_1_81_Update/ca
      -- 
    ca_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1_81_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_sample_start_
      -- 
    inputPort_1_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(12);
      gj_inputPort_1_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(60) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(66);
      gj_inputPort_1_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_sample_start__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(39) <= inputPort_1_Daemon_CP_3_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_update_start__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(41) <= inputPort_1_Daemon_CP_3_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_update_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_loopback_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(43) <= inputPort_1_Daemon_CP_3_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_loopback_sample_req_ps
      -- 
    phi_stmt_82_loopback_sample_req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_82_loopback_sample_req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(44), ack => phi_stmt_82_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_entry_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(45) <= inputPort_1_Daemon_CP_3_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_entry_sample_req_ps
      -- 
    phi_stmt_82_entry_sample_req_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_82_entry_sample_req_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(46), ack => phi_stmt_82_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/phi_stmt_82_phi_mux_ack_ps
      -- 
    phi_stmt_82_phi_mux_ack_110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_82_ack_0, ack => inputPort_1_Daemon_CP_3_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/konst_84_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/konst_84_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/konst_84_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/konst_84_sample_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/konst_84_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/konst_84_update_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/konst_84_update_completed__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(50) <= inputPort_1_Daemon_CP_3_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/konst_84_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(49), ack => inputPort_1_Daemon_CP_3_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_Sample/req
      -- 
    req_131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(52), ack => next_last_dest_id_117_85_buf_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_update_start_
      -- CP-element group 53: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_Update/req
      -- 
    req_136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(53), ack => next_last_dest_id_117_85_buf_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_Sample/ack
      -- 
    ack_132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_117_85_buf_ack_0, ack => inputPort_1_Daemon_CP_3_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/R_next_last_dest_id_85_Update/ack
      -- 
    ack_137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_117_85_buf_ack_1, ack => inputPort_1_Daemon_CP_3_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_Sample/req
      -- 
    req_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(56), ack => WPIPE_noblock_obuf_1_1_129_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(58);
      gj_inputPort_1_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_update_start_
      -- CP-element group 57: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_Update/req
      -- 
    ack_147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_1_129_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(57)); -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(57), ack => WPIPE_noblock_obuf_1_1_129_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_1_129_Update/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_1_129_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_Sample/req
      -- 
    req_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(59), ack => WPIPE_noblock_obuf_1_2_138_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(61);
      gj_inputPort_1_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_update_start_
      -- CP-element group 60: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_Update/req
      -- 
    ack_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_2_138_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(60)); -- 
    req_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(60), ack => WPIPE_noblock_obuf_1_2_138_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_2_138_Update/ack
      -- 
    ack_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_2_138_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_Sample/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(62), ack => WPIPE_noblock_obuf_1_3_147_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(64);
      gj_inputPort_1_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_update_start_
      -- CP-element group 63: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_Update/req
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_3_147_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(63)); -- 
    req_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(63), ack => WPIPE_noblock_obuf_1_3_147_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_3_147_Update/ack
      -- 
    ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_3_147_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_Sample/req
      -- 
    req_188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(65), ack => WPIPE_noblock_obuf_1_4_156_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(67);
      gj_inputPort_1_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_update_start_
      -- CP-element group 66: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_Update/req
      -- 
    ack_189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_4_156_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(66)); -- 
    req_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(66), ack => WPIPE_noblock_obuf_1_4_156_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/WPIPE_noblock_obuf_1_4_156_Update/ack
      -- 
    ack_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_4_156_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(9), ack => inputPort_1_Daemon_CP_3_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_71/do_while_stmt_72/do_while_stmt_72_loop_body/$exit
      -- 
    inputPort_1_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(12) & inputPort_1_Daemon_CP_3_elements(58) & inputPort_1_Daemon_CP_3_elements(61) & inputPort_1_Daemon_CP_3_elements(64) & inputPort_1_Daemon_CP_3_elements(67);
      gj_inputPort_1_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_71/do_while_stmt_72/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_71/do_while_stmt_72/loop_exit/ack
      -- 
    ack_199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_72_branch_ack_0, ack => inputPort_1_Daemon_CP_3_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_71/do_while_stmt_72/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_71/do_while_stmt_72/loop_taken/ack
      -- 
    ack_203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_72_branch_ack_1, ack => inputPort_1_Daemon_CP_3_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_71/do_while_stmt_72/$exit
      -- 
    inputPort_1_Daemon_CP_3_elements(72) <= inputPort_1_Daemon_CP_3_elements(3);
    inputPort_1_Daemon_do_while_stmt_72_terminator_204: loop_terminator -- 
      generic map (name => " inputPort_1_Daemon_do_while_stmt_72_terminator_204", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_1_Daemon_CP_3_elements(6),loop_continue => inputPort_1_Daemon_CP_3_elements(71),loop_terminate => inputPort_1_Daemon_CP_3_elements(70),loop_back => inputPort_1_Daemon_CP_3_elements(4),loop_exit => inputPort_1_Daemon_CP_3_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_74_phi_seq_76_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_1_Daemon_CP_3_elements(19);
      inputPort_1_Daemon_CP_3_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_1_Daemon_CP_3_elements(26);
      inputPort_1_Daemon_CP_3_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_1_Daemon_CP_3_elements(27);
      inputPort_1_Daemon_CP_3_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_1_Daemon_CP_3_elements(21);
      inputPort_1_Daemon_CP_3_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_1_Daemon_CP_3_elements(28);
      inputPort_1_Daemon_CP_3_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_1_Daemon_CP_3_elements(30);
      inputPort_1_Daemon_CP_3_elements(22) <= phi_mux_reqs(1);
      phi_stmt_74_phi_seq_76 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_74_phi_seq_76") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_1_Daemon_CP_3_elements(11), 
          phi_sample_ack => inputPort_1_Daemon_CP_3_elements(17), 
          phi_update_req => inputPort_1_Daemon_CP_3_elements(13), 
          phi_update_ack => inputPort_1_Daemon_CP_3_elements(18), 
          phi_mux_ack => inputPort_1_Daemon_CP_3_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_82_phi_seq_138_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_1_Daemon_CP_3_elements(45);
      inputPort_1_Daemon_CP_3_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_1_Daemon_CP_3_elements(48);
      inputPort_1_Daemon_CP_3_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_1_Daemon_CP_3_elements(50);
      inputPort_1_Daemon_CP_3_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_1_Daemon_CP_3_elements(43);
      inputPort_1_Daemon_CP_3_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_1_Daemon_CP_3_elements(54);
      inputPort_1_Daemon_CP_3_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_1_Daemon_CP_3_elements(55);
      inputPort_1_Daemon_CP_3_elements(44) <= phi_mux_reqs(1);
      phi_stmt_82_phi_seq_138 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_82_phi_seq_138") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_1_Daemon_CP_3_elements(39), 
          phi_sample_ack => inputPort_1_Daemon_CP_3_elements(40), 
          phi_update_req => inputPort_1_Daemon_CP_3_elements(41), 
          phi_update_ack => inputPort_1_Daemon_CP_3_elements(42), 
          phi_mux_ack => inputPort_1_Daemon_CP_3_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_28_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_1_Daemon_CP_3_elements(7);
        preds(1)  <= inputPort_1_Daemon_CP_3_elements(8);
        entry_tmerge_28 : transition_merge -- 
          generic map(name => " entry_tmerge_28")
          port map (preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_1_81_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_119_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_106_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_109_wire : std_logic_vector(15 downto 0);
    signal count_down_74 : std_logic_vector(15 downto 0);
    signal data_to_outport_122 : std_logic_vector(32 downto 0);
    signal dest_id_97 : std_logic_vector(7 downto 0);
    signal input_word_79 : std_logic_vector(31 downto 0);
    signal konst_105_wire_constant : std_logic_vector(15 downto 0);
    signal konst_108_wire_constant : std_logic_vector(15 downto 0);
    signal konst_125_wire_constant : std_logic_vector(7 downto 0);
    signal konst_134_wire_constant : std_logic_vector(7 downto 0);
    signal konst_143_wire_constant : std_logic_vector(7 downto 0);
    signal konst_152_wire_constant : std_logic_vector(7 downto 0);
    signal konst_170_wire_constant : std_logic_vector(0 downto 0);
    signal konst_84_wire_constant : std_logic_vector(7 downto 0);
    signal konst_89_wire_constant : std_logic_vector(15 downto 0);
    signal last_dest_id_82 : std_logic_vector(7 downto 0);
    signal new_packet_91 : std_logic_vector(0 downto 0);
    signal next_count_down_111 : std_logic_vector(15 downto 0);
    signal next_count_down_111_76_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_117 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_117_85_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_101 : std_logic_vector(15 downto 0);
    signal send_to_1_127 : std_logic_vector(0 downto 0);
    signal send_to_2_136 : std_logic_vector(0 downto 0);
    signal send_to_3_145 : std_logic_vector(0 downto 0);
    signal send_to_4_154 : std_logic_vector(0 downto 0);
    signal type_cast_78_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_119_wire_constant <= "1";
    konst_105_wire_constant <= "0000000000000001";
    konst_108_wire_constant <= "0000000000000001";
    konst_125_wire_constant <= "00000001";
    konst_134_wire_constant <= "00000010";
    konst_143_wire_constant <= "00000011";
    konst_152_wire_constant <= "00000100";
    konst_170_wire_constant <= "1";
    konst_84_wire_constant <= "00000000";
    konst_89_wire_constant <= "0000000000000000";
    type_cast_78_wire_constant <= "0000000000000000";
    phi_stmt_74: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_count_down_111_76_buffered & type_cast_78_wire_constant;
      req <= phi_stmt_74_req_0 & phi_stmt_74_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_74",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_74_ack_0,
          idata => idata,
          odata => count_down_74,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_74
    phi_stmt_82: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_84_wire_constant & next_last_dest_id_117_85_buffered;
      req <= phi_stmt_82_req_0 & phi_stmt_82_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_82",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_82_ack_0,
          idata => idata,
          odata => last_dest_id_82,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_82
    -- flow-through select operator MUX_110_inst
    next_count_down_111 <= SUB_u16_u16_106_wire when (new_packet_91(0) /=  '0') else SUB_u16_u16_109_wire;
    -- flow-through select operator MUX_116_inst
    next_last_dest_id_117 <= dest_id_97 when (new_packet_91(0) /=  '0') else last_dest_id_82;
    -- flow-through slice operator slice_100_inst
    pkt_length_101 <= input_word_79(23 downto 8);
    -- flow-through slice operator slice_96_inst
    dest_id_97 <= input_word_79(31 downto 24);
    next_count_down_111_76_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_111_76_buf_req_0;
      next_count_down_111_76_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_111_76_buf_req_1;
      next_count_down_111_76_buf_ack_1<= rack(0);
      next_count_down_111_76_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_111_76_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_111_76_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_117_85_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_117_85_buf_req_0;
      next_last_dest_id_117_85_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_117_85_buf_req_1;
      next_last_dest_id_117_85_buf_ack_1<= rack(0);
      next_last_dest_id_117_85_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_117_85_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_117_85_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_79
    process(RPIPE_in_data_1_81_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_1_81_wire(31 downto 0);
      input_word_79 <= tmp_var; -- 
    end process;
    do_while_stmt_72_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_170_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_72_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_72_branch_req_0,
          ack0 => do_while_stmt_72_branch_ack_0,
          ack1 => do_while_stmt_72_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_121_inst
    process(R_ONE_1_119_wire_constant, input_word_79) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_119_wire_constant, input_word_79, tmp_var);
      data_to_outport_122 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_90_inst
    process(count_down_74) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_74, konst_89_wire_constant, tmp_var);
      new_packet_91 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_126_inst
    process(next_last_dest_id_117) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_117, konst_125_wire_constant, tmp_var);
      send_to_1_127 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_135_inst
    process(next_last_dest_id_117) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_117, konst_134_wire_constant, tmp_var);
      send_to_2_136 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_144_inst
    process(next_last_dest_id_117) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_117, konst_143_wire_constant, tmp_var);
      send_to_3_145 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_153_inst
    process(next_last_dest_id_117) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_117, konst_152_wire_constant, tmp_var);
      send_to_4_154 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_106_inst
    process(pkt_length_101) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_101, konst_105_wire_constant, tmp_var);
      SUB_u16_u16_106_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_109_inst
    process(count_down_74) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_74, konst_108_wire_constant, tmp_var);
      SUB_u16_u16_109_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_1_81_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_1_81_inst_req_0;
      RPIPE_in_data_1_81_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_1_81_inst_req_1;
      RPIPE_in_data_1_81_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_1_81_wire <= data_out(31 downto 0);
      in_data_1_read_0_gI: SplitGuardInterface generic map(name => "in_data_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_1_read_0: InputPortRevised -- 
        generic map ( name => "in_data_1_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_1_pipe_read_req(0),
          oack => in_data_1_pipe_read_ack(0),
          odata => in_data_1_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_1_1_129_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_1_129_inst_req_0;
      WPIPE_noblock_obuf_1_1_129_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_1_129_inst_req_1;
      WPIPE_noblock_obuf_1_1_129_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_127(0);
      data_in <= data_to_outport_122;
      noblock_obuf_1_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_1_pipe_write_req(0),
          oack => noblock_obuf_1_1_pipe_write_ack(0),
          odata => noblock_obuf_1_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_1_2_138_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_2_138_inst_req_0;
      WPIPE_noblock_obuf_1_2_138_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_2_138_inst_req_1;
      WPIPE_noblock_obuf_1_2_138_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_136(0);
      data_in <= data_to_outport_122;
      noblock_obuf_1_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_2_pipe_write_req(0),
          oack => noblock_obuf_1_2_pipe_write_ack(0),
          odata => noblock_obuf_1_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_1_3_147_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_3_147_inst_req_0;
      WPIPE_noblock_obuf_1_3_147_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_3_147_inst_req_1;
      WPIPE_noblock_obuf_1_3_147_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_145(0);
      data_in <= data_to_outport_122;
      noblock_obuf_1_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_3_pipe_write_req(0),
          oack => noblock_obuf_1_3_pipe_write_ack(0),
          odata => noblock_obuf_1_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_1_4_156_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_4_156_inst_req_0;
      WPIPE_noblock_obuf_1_4_156_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_4_156_inst_req_1;
      WPIPE_noblock_obuf_1_4_156_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_154(0);
      data_in <= data_to_outport_122;
      noblock_obuf_1_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_4_pipe_write_req(0),
          oack => noblock_obuf_1_4_pipe_write_ack(0),
          odata => noblock_obuf_1_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_1_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_2_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_2_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_2_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_2_Daemon;
architecture inputPort_2_Daemon_arch of inputPort_2_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_2_Daemon_CP_205_start: Boolean;
  signal inputPort_2_Daemon_CP_205_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_noblock_obuf_2_3_250_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_250_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_250_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_3_250_inst_ack_1 : boolean;
  signal do_while_stmt_175_branch_req_0 : boolean;
  signal phi_stmt_177_req_1 : boolean;
  signal phi_stmt_177_req_0 : boolean;
  signal phi_stmt_177_ack_0 : boolean;
  signal next_count_down_214_181_buf_req_0 : boolean;
  signal next_count_down_214_181_buf_ack_0 : boolean;
  signal next_count_down_214_181_buf_req_1 : boolean;
  signal next_count_down_214_181_buf_ack_1 : boolean;
  signal RPIPE_in_data_2_184_inst_req_0 : boolean;
  signal RPIPE_in_data_2_184_inst_ack_0 : boolean;
  signal RPIPE_in_data_2_184_inst_req_1 : boolean;
  signal RPIPE_in_data_2_184_inst_ack_1 : boolean;
  signal phi_stmt_185_req_0 : boolean;
  signal phi_stmt_185_req_1 : boolean;
  signal phi_stmt_185_ack_0 : boolean;
  signal next_last_dest_id_220_187_buf_req_0 : boolean;
  signal next_last_dest_id_220_187_buf_ack_0 : boolean;
  signal next_last_dest_id_220_187_buf_req_1 : boolean;
  signal next_last_dest_id_220_187_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_1_232_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_1_232_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_1_232_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_1_232_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_241_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_2_241_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_2_241_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_241_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_259_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_4_259_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_4_259_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_259_inst_ack_1 : boolean;
  signal do_while_stmt_175_branch_ack_0 : boolean;
  signal do_while_stmt_175_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_2_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_2_Daemon_CP_205_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_2_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_2_Daemon_CP_205: Block -- control-path 
    signal inputPort_2_Daemon_CP_205_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_2_Daemon_CP_205_elements(0) <= inputPort_2_Daemon_CP_205_start;
    inputPort_2_Daemon_CP_205_symbol <= inputPort_2_Daemon_CP_205_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_174/$entry
      -- CP-element group 0: 	 branch_block_stmt_174/branch_block_stmt_174__entry__
      -- CP-element group 0: 	 branch_block_stmt_174/do_while_stmt_175__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_174/$exit
      -- CP-element group 1: 	 branch_block_stmt_174/branch_block_stmt_174__exit__
      -- CP-element group 1: 	 branch_block_stmt_174/do_while_stmt_175__exit__
      -- 
    inputPort_2_Daemon_CP_205_elements(1) <= inputPort_2_Daemon_CP_205_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_174/do_while_stmt_175/$entry
      -- CP-element group 2: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175__entry__
      -- 
    inputPort_2_Daemon_CP_205_elements(2) <= inputPort_2_Daemon_CP_205_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175__exit__
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_174/do_while_stmt_175/loop_back
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	70 
    -- CP-element group 5: 	71 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_174/do_while_stmt_175/condition_done
      -- CP-element group 5: 	 branch_block_stmt_174/do_while_stmt_175/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_174/do_while_stmt_175/loop_taken/$entry
      -- 
    inputPort_2_Daemon_CP_205_elements(5) <= inputPort_2_Daemon_CP_205_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_174/do_while_stmt_175/loop_body_done
      -- 
    inputPort_2_Daemon_CP_205_elements(6) <= inputPort_2_Daemon_CP_205_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/back_edge_to_loop_body
      -- 
    inputPort_2_Daemon_CP_205_elements(7) <= inputPort_2_Daemon_CP_205_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/first_time_through_loop_body
      -- 
    inputPort_2_Daemon_CP_205_elements(8) <= inputPort_2_Daemon_CP_205_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	68 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_182_sample_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/condition_evaluated
      -- 
    condition_evaluated_229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(10), ack => do_while_stmt_175_branch_req_0); -- 
    inputPort_2_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(14) & inputPort_2_Daemon_CP_205_elements(68);
      gj_inputPort_2_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_sample_start__ps
      -- 
    inputPort_2_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(15) & inputPort_2_Daemon_CP_205_elements(37) & inputPort_2_Daemon_CP_205_elements(14);
      gj_inputPort_2_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_182_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_sample_completed_
      -- 
    inputPort_2_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(17) & inputPort_2_Daemon_CP_205_elements(35) & inputPort_2_Daemon_CP_205_elements(40);
      gj_inputPort_2_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_update_start__ps
      -- 
    inputPort_2_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(16) & inputPort_2_Daemon_CP_205_elements(32) & inputPort_2_Daemon_CP_205_elements(38);
      gj_inputPort_2_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_2_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42);
      gj_inputPort_2_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_sample_start_
      -- 
    inputPort_2_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_sample_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_update_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_loopback_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(19) <= inputPort_2_Daemon_CP_205_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_loopback_sample_req_ps
      -- 
    phi_stmt_177_loopback_sample_req_244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_177_loopback_sample_req_244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(20), ack => phi_stmt_177_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_entry_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(21) <= inputPort_2_Daemon_CP_205_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_entry_sample_req_ps
      -- 
    phi_stmt_177_entry_sample_req_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_177_entry_sample_req_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(22), ack => phi_stmt_177_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_177_phi_mux_ack_ps
      -- 
    phi_stmt_177_phi_mux_ack_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_177_ack_0, ack => inputPort_2_Daemon_CP_205_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/type_cast_180_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/type_cast_180_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/type_cast_180_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/type_cast_180_sample_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/type_cast_180_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/type_cast_180_update_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/type_cast_180_update_completed__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(26) <= inputPort_2_Daemon_CP_205_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/type_cast_180_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(25), ack => inputPort_2_Daemon_CP_205_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_Sample/req
      -- 
    req_271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(28), ack => next_count_down_214_181_buf_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_update_start_
      -- CP-element group 29: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_Update/req
      -- 
    req_276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(29), ack => next_count_down_214_181_buf_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_Sample/ack
      -- 
    ack_272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_214_181_buf_ack_0, ack => inputPort_2_Daemon_CP_205_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_count_down_181_Update/ack
      -- 
    ack_277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_214_181_buf_ack_1, ack => inputPort_2_Daemon_CP_205_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_182_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_Sample/rr
      -- 
    rr_290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(33), ack => RPIPE_in_data_2_184_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(11) & inputPort_2_Daemon_CP_205_elements(36);
      gj_inputPort_2_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_update_start_
      -- CP-element group 34: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_Update/cr
      -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(34), ack => RPIPE_in_data_2_184_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(13) & inputPort_2_Daemon_CP_205_elements(35);
      gj_inputPort_2_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_Sample/ra
      -- 
    ra_291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2_184_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_182_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/RPIPE_in_data_2_184_Update/ca
      -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2_184_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_sample_start_
      -- 
    inputPort_2_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_sample_start__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(39) <= inputPort_2_Daemon_CP_205_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_sample_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_update_start__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(41) <= inputPort_2_Daemon_CP_205_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_update_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_loopback_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(43) <= inputPort_2_Daemon_CP_205_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_loopback_sample_req_ps
      -- 
    phi_stmt_185_loopback_sample_req_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_185_loopback_sample_req_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(44), ack => phi_stmt_185_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_entry_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(45) <= inputPort_2_Daemon_CP_205_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_entry_sample_req_ps
      -- 
    phi_stmt_185_entry_sample_req_309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_185_entry_sample_req_309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(46), ack => phi_stmt_185_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/phi_stmt_185_phi_mux_ack_ps
      -- 
    phi_stmt_185_phi_mux_ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_185_ack_0, ack => inputPort_2_Daemon_CP_205_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_Sample/req
      -- 
    req_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(48), ack => next_last_dest_id_220_187_buf_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_update_start_
      -- CP-element group 49: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_Update/req
      -- 
    req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(49), ack => next_last_dest_id_220_187_buf_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_sample_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_Sample/ack
      -- 
    ack_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_220_187_buf_ack_0, ack => inputPort_2_Daemon_CP_205_elements(50)); -- 
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_update_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/R_next_last_dest_id_187_Update/ack
      -- 
    ack_331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_220_187_buf_ack_1, ack => inputPort_2_Daemon_CP_205_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/konst_188_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/konst_188_sample_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/konst_188_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/konst_188_sample_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/konst_188_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/konst_188_update_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/konst_188_update_completed__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(54) <= inputPort_2_Daemon_CP_205_elements(55);
    -- CP-element group 55:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	54 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/konst_188_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(55) is a control-delay.
    cp_element_55_delay: control_delay_element  generic map(name => " 55_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(53), ack => inputPort_2_Daemon_CP_205_elements(55), clk => clk, reset =>reset);
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_Sample/req
      -- 
    req_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(56), ack => WPIPE_noblock_obuf_2_1_232_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(58);
      gj_inputPort_2_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_update_start_
      -- CP-element group 57: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_Update/req
      -- 
    ack_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_1_232_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(57)); -- 
    req_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(57), ack => WPIPE_noblock_obuf_2_1_232_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_1_232_Update/ack
      -- 
    ack_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_1_232_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_Sample/req
      -- 
    req_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(59), ack => WPIPE_noblock_obuf_2_2_241_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(61);
      gj_inputPort_2_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_update_start_
      -- CP-element group 60: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_Update/req
      -- 
    ack_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_2_241_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(60)); -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(60), ack => WPIPE_noblock_obuf_2_2_241_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_2_241_Update/ack
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_2_241_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_sample_start_
      -- 
    req_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(62), ack => WPIPE_noblock_obuf_2_3_250_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(64);
      gj_inputPort_2_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_update_start_
      -- CP-element group 63: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_Update/req
      -- CP-element group 63: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_sample_completed_
      -- 
    ack_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_3_250_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(63)); -- 
    req_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(63), ack => WPIPE_noblock_obuf_2_3_250_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_3_250_Update/ack
      -- 
    ack_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_3_250_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_Sample/req
      -- 
    req_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(65), ack => WPIPE_noblock_obuf_2_4_259_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(67);
      gj_inputPort_2_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_update_start_
      -- CP-element group 66: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_Update/req
      -- 
    ack_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_4_259_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(66)); -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(66), ack => WPIPE_noblock_obuf_2_4_259_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/WPIPE_noblock_obuf_2_4_259_Update/ack
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_4_259_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(9), ack => inputPort_2_Daemon_CP_205_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_174/do_while_stmt_175/do_while_stmt_175_loop_body/$exit
      -- 
    inputPort_2_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(12) & inputPort_2_Daemon_CP_205_elements(58) & inputPort_2_Daemon_CP_205_elements(61) & inputPort_2_Daemon_CP_205_elements(64) & inputPort_2_Daemon_CP_205_elements(67);
      gj_inputPort_2_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_174/do_while_stmt_175/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_174/do_while_stmt_175/loop_exit/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_175_branch_ack_0, ack => inputPort_2_Daemon_CP_205_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_174/do_while_stmt_175/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_174/do_while_stmt_175/loop_taken/ack
      -- 
    ack_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_175_branch_ack_1, ack => inputPort_2_Daemon_CP_205_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_174/do_while_stmt_175/$exit
      -- 
    inputPort_2_Daemon_CP_205_elements(72) <= inputPort_2_Daemon_CP_205_elements(3);
    inputPort_2_Daemon_do_while_stmt_175_terminator_406: loop_terminator -- 
      generic map (name => " inputPort_2_Daemon_do_while_stmt_175_terminator_406", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_2_Daemon_CP_205_elements(6),loop_continue => inputPort_2_Daemon_CP_205_elements(71),loop_terminate => inputPort_2_Daemon_CP_205_elements(70),loop_back => inputPort_2_Daemon_CP_205_elements(4),loop_exit => inputPort_2_Daemon_CP_205_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_177_phi_seq_278_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_2_Daemon_CP_205_elements(21);
      inputPort_2_Daemon_CP_205_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_2_Daemon_CP_205_elements(24);
      inputPort_2_Daemon_CP_205_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_2_Daemon_CP_205_elements(26);
      inputPort_2_Daemon_CP_205_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_2_Daemon_CP_205_elements(19);
      inputPort_2_Daemon_CP_205_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_2_Daemon_CP_205_elements(30);
      inputPort_2_Daemon_CP_205_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_2_Daemon_CP_205_elements(31);
      inputPort_2_Daemon_CP_205_elements(20) <= phi_mux_reqs(1);
      phi_stmt_177_phi_seq_278 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_177_phi_seq_278") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_2_Daemon_CP_205_elements(11), 
          phi_sample_ack => inputPort_2_Daemon_CP_205_elements(17), 
          phi_update_req => inputPort_2_Daemon_CP_205_elements(13), 
          phi_update_ack => inputPort_2_Daemon_CP_205_elements(18), 
          phi_mux_ack => inputPort_2_Daemon_CP_205_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_185_phi_seq_340_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_2_Daemon_CP_205_elements(43);
      inputPort_2_Daemon_CP_205_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_2_Daemon_CP_205_elements(50);
      inputPort_2_Daemon_CP_205_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_2_Daemon_CP_205_elements(51);
      inputPort_2_Daemon_CP_205_elements(44) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_2_Daemon_CP_205_elements(45);
      inputPort_2_Daemon_CP_205_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_2_Daemon_CP_205_elements(52);
      inputPort_2_Daemon_CP_205_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_2_Daemon_CP_205_elements(54);
      inputPort_2_Daemon_CP_205_elements(46) <= phi_mux_reqs(1);
      phi_stmt_185_phi_seq_340 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_185_phi_seq_340") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_2_Daemon_CP_205_elements(39), 
          phi_sample_ack => inputPort_2_Daemon_CP_205_elements(40), 
          phi_update_req => inputPort_2_Daemon_CP_205_elements(41), 
          phi_update_ack => inputPort_2_Daemon_CP_205_elements(42), 
          phi_mux_ack => inputPort_2_Daemon_CP_205_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_230_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_2_Daemon_CP_205_elements(7);
        preds(1)  <= inputPort_2_Daemon_CP_205_elements(8);
        entry_tmerge_230 : transition_merge -- 
          generic map(name => " entry_tmerge_230")
          port map (preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_2_184_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_222_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_209_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_212_wire : std_logic_vector(15 downto 0);
    signal count_down_177 : std_logic_vector(15 downto 0);
    signal data_to_outport_225 : std_logic_vector(32 downto 0);
    signal dest_id_200 : std_logic_vector(7 downto 0);
    signal input_word_182 : std_logic_vector(31 downto 0);
    signal konst_188_wire_constant : std_logic_vector(7 downto 0);
    signal konst_192_wire_constant : std_logic_vector(15 downto 0);
    signal konst_208_wire_constant : std_logic_vector(15 downto 0);
    signal konst_211_wire_constant : std_logic_vector(15 downto 0);
    signal konst_228_wire_constant : std_logic_vector(7 downto 0);
    signal konst_237_wire_constant : std_logic_vector(7 downto 0);
    signal konst_246_wire_constant : std_logic_vector(7 downto 0);
    signal konst_255_wire_constant : std_logic_vector(7 downto 0);
    signal konst_273_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_185 : std_logic_vector(7 downto 0);
    signal new_packet_194 : std_logic_vector(0 downto 0);
    signal next_count_down_214 : std_logic_vector(15 downto 0);
    signal next_count_down_214_181_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_220 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_220_187_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_204 : std_logic_vector(15 downto 0);
    signal send_to_1_230 : std_logic_vector(0 downto 0);
    signal send_to_2_239 : std_logic_vector(0 downto 0);
    signal send_to_3_248 : std_logic_vector(0 downto 0);
    signal send_to_4_257 : std_logic_vector(0 downto 0);
    signal type_cast_180_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_222_wire_constant <= "1";
    konst_188_wire_constant <= "00000000";
    konst_192_wire_constant <= "0000000000000000";
    konst_208_wire_constant <= "0000000000000001";
    konst_211_wire_constant <= "0000000000000001";
    konst_228_wire_constant <= "00000001";
    konst_237_wire_constant <= "00000010";
    konst_246_wire_constant <= "00000011";
    konst_255_wire_constant <= "00000100";
    konst_273_wire_constant <= "1";
    type_cast_180_wire_constant <= "0000000000000000";
    phi_stmt_177: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_180_wire_constant & next_count_down_214_181_buffered;
      req <= phi_stmt_177_req_0 & phi_stmt_177_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_177",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_177_ack_0,
          idata => idata,
          odata => count_down_177,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_177
    phi_stmt_185: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_last_dest_id_220_187_buffered & konst_188_wire_constant;
      req <= phi_stmt_185_req_0 & phi_stmt_185_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_185",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_185_ack_0,
          idata => idata,
          odata => last_dest_id_185,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_185
    -- flow-through select operator MUX_213_inst
    next_count_down_214 <= SUB_u16_u16_209_wire when (new_packet_194(0) /=  '0') else SUB_u16_u16_212_wire;
    -- flow-through select operator MUX_219_inst
    next_last_dest_id_220 <= dest_id_200 when (new_packet_194(0) /=  '0') else last_dest_id_185;
    -- flow-through slice operator slice_199_inst
    dest_id_200 <= input_word_182(31 downto 24);
    -- flow-through slice operator slice_203_inst
    pkt_length_204 <= input_word_182(23 downto 8);
    next_count_down_214_181_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_214_181_buf_req_0;
      next_count_down_214_181_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_214_181_buf_req_1;
      next_count_down_214_181_buf_ack_1<= rack(0);
      next_count_down_214_181_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_214_181_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_214_181_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_220_187_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_220_187_buf_req_0;
      next_last_dest_id_220_187_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_220_187_buf_req_1;
      next_last_dest_id_220_187_buf_ack_1<= rack(0);
      next_last_dest_id_220_187_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_220_187_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_220_187_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_182
    process(RPIPE_in_data_2_184_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_2_184_wire(31 downto 0);
      input_word_182 <= tmp_var; -- 
    end process;
    do_while_stmt_175_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_273_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_175_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_175_branch_req_0,
          ack0 => do_while_stmt_175_branch_ack_0,
          ack1 => do_while_stmt_175_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_224_inst
    process(R_ONE_1_222_wire_constant, input_word_182) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_222_wire_constant, input_word_182, tmp_var);
      data_to_outport_225 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_193_inst
    process(count_down_177) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_177, konst_192_wire_constant, tmp_var);
      new_packet_194 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_229_inst
    process(next_last_dest_id_220) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_220, konst_228_wire_constant, tmp_var);
      send_to_1_230 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_238_inst
    process(next_last_dest_id_220) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_220, konst_237_wire_constant, tmp_var);
      send_to_2_239 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_247_inst
    process(next_last_dest_id_220) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_220, konst_246_wire_constant, tmp_var);
      send_to_3_248 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_256_inst
    process(next_last_dest_id_220) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_220, konst_255_wire_constant, tmp_var);
      send_to_4_257 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_209_inst
    process(pkt_length_204) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_204, konst_208_wire_constant, tmp_var);
      SUB_u16_u16_209_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_212_inst
    process(count_down_177) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_177, konst_211_wire_constant, tmp_var);
      SUB_u16_u16_212_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_2_184_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_2_184_inst_req_0;
      RPIPE_in_data_2_184_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_2_184_inst_req_1;
      RPIPE_in_data_2_184_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_2_184_wire <= data_out(31 downto 0);
      in_data_2_read_0_gI: SplitGuardInterface generic map(name => "in_data_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_2_read_0: InputPortRevised -- 
        generic map ( name => "in_data_2_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_2_pipe_read_req(0),
          oack => in_data_2_pipe_read_ack(0),
          odata => in_data_2_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_2_1_232_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_1_232_inst_req_0;
      WPIPE_noblock_obuf_2_1_232_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_1_232_inst_req_1;
      WPIPE_noblock_obuf_2_1_232_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_230(0);
      data_in <= data_to_outport_225;
      noblock_obuf_2_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_1_pipe_write_req(0),
          oack => noblock_obuf_2_1_pipe_write_ack(0),
          odata => noblock_obuf_2_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_2_2_241_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_2_241_inst_req_0;
      WPIPE_noblock_obuf_2_2_241_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_2_241_inst_req_1;
      WPIPE_noblock_obuf_2_2_241_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_239(0);
      data_in <= data_to_outport_225;
      noblock_obuf_2_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_2_pipe_write_req(0),
          oack => noblock_obuf_2_2_pipe_write_ack(0),
          odata => noblock_obuf_2_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_2_3_250_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_3_250_inst_req_0;
      WPIPE_noblock_obuf_2_3_250_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_3_250_inst_req_1;
      WPIPE_noblock_obuf_2_3_250_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_248(0);
      data_in <= data_to_outport_225;
      noblock_obuf_2_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_3_pipe_write_req(0),
          oack => noblock_obuf_2_3_pipe_write_ack(0),
          odata => noblock_obuf_2_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_2_4_259_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_4_259_inst_req_0;
      WPIPE_noblock_obuf_2_4_259_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_4_259_inst_req_1;
      WPIPE_noblock_obuf_2_4_259_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_257(0);
      data_in <= data_to_outport_225;
      noblock_obuf_2_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_4_pipe_write_req(0),
          oack => noblock_obuf_2_4_pipe_write_ack(0),
          odata => noblock_obuf_2_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_2_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_3_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_3_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_3_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_3_Daemon;
architecture inputPort_3_Daemon_arch of inputPort_3_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_3_Daemon_CP_407_start: Boolean;
  signal inputPort_3_Daemon_CP_407_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal next_last_dest_id_323_291_buf_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_4_362_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_362_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_353_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_1_335_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_344_inst_ack_1 : boolean;
  signal next_count_down_317_284_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_353_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_344_inst_req_1 : boolean;
  signal phi_stmt_288_ack_0 : boolean;
  signal RPIPE_in_data_3_287_inst_ack_1 : boolean;
  signal next_count_down_317_284_buf_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_1_335_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_1_335_inst_req_1 : boolean;
  signal do_while_stmt_278_branch_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_2_344_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_344_inst_req_0 : boolean;
  signal next_last_dest_id_323_291_buf_req_0 : boolean;
  signal RPIPE_in_data_3_287_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_1_335_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_4_362_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_4_362_inst_req_0 : boolean;
  signal next_count_down_317_284_buf_ack_0 : boolean;
  signal do_while_stmt_278_branch_ack_0 : boolean;
  signal next_count_down_317_284_buf_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_3_353_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_353_inst_req_1 : boolean;
  signal phi_stmt_288_req_0 : boolean;
  signal phi_stmt_288_req_1 : boolean;
  signal RPIPE_in_data_3_287_inst_ack_0 : boolean;
  signal RPIPE_in_data_3_287_inst_req_0 : boolean;
  signal next_last_dest_id_323_291_buf_ack_1 : boolean;
  signal next_last_dest_id_323_291_buf_req_1 : boolean;
  signal phi_stmt_280_ack_0 : boolean;
  signal phi_stmt_280_req_0 : boolean;
  signal phi_stmt_280_req_1 : boolean;
  signal do_while_stmt_278_branch_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_3_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_3_Daemon_CP_407_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_3_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_3_Daemon_CP_407: Block -- control-path 
    signal inputPort_3_Daemon_CP_407_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_3_Daemon_CP_407_elements(0) <= inputPort_3_Daemon_CP_407_start;
    inputPort_3_Daemon_CP_407_symbol <= inputPort_3_Daemon_CP_407_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_277/$entry
      -- CP-element group 0: 	 branch_block_stmt_277/branch_block_stmt_277__entry__
      -- CP-element group 0: 	 branch_block_stmt_277/do_while_stmt_278__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_277/$exit
      -- CP-element group 1: 	 branch_block_stmt_277/branch_block_stmt_277__exit__
      -- CP-element group 1: 	 branch_block_stmt_277/do_while_stmt_278__exit__
      -- 
    inputPort_3_Daemon_CP_407_elements(1) <= inputPort_3_Daemon_CP_407_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_277/do_while_stmt_278/$entry
      -- CP-element group 2: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278__entry__
      -- 
    inputPort_3_Daemon_CP_407_elements(2) <= inputPort_3_Daemon_CP_407_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278__exit__
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_277/do_while_stmt_278/loop_back
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	70 
    -- CP-element group 5: 	71 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_277/do_while_stmt_278/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_277/do_while_stmt_278/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_277/do_while_stmt_278/condition_done
      -- 
    inputPort_3_Daemon_CP_407_elements(5) <= inputPort_3_Daemon_CP_407_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_277/do_while_stmt_278/loop_body_done
      -- 
    inputPort_3_Daemon_CP_407_elements(6) <= inputPort_3_Daemon_CP_407_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/back_edge_to_loop_body
      -- 
    inputPort_3_Daemon_CP_407_elements(7) <= inputPort_3_Daemon_CP_407_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/first_time_through_loop_body
      -- 
    inputPort_3_Daemon_CP_407_elements(8) <= inputPort_3_Daemon_CP_407_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	68 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_285_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/loop_body_start
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	68 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/condition_evaluated
      -- 
    condition_evaluated_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(10), ack => do_while_stmt_278_branch_req_0); -- 
    inputPort_3_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(68) & inputPort_3_Daemon_CP_407_elements(14);
      gj_inputPort_3_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/aggregated_phi_sample_req
      -- 
    inputPort_3_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(15) & inputPort_3_Daemon_CP_407_elements(37) & inputPort_3_Daemon_CP_407_elements(14);
      gj_inputPort_3_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_285_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_sample_completed_
      -- 
    inputPort_3_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(17) & inputPort_3_Daemon_CP_407_elements(35) & inputPort_3_Daemon_CP_407_elements(40);
      gj_inputPort_3_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_update_start__ps
      -- 
    inputPort_3_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(16) & inputPort_3_Daemon_CP_407_elements(32) & inputPort_3_Daemon_CP_407_elements(38);
      gj_inputPort_3_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_3_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42);
      gj_inputPort_3_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_sample_start_
      -- 
    inputPort_3_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(12);
      gj_inputPort_3_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_sample_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_loopback_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(19) <= inputPort_3_Daemon_CP_407_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_loopback_sample_req
      -- 
    phi_stmt_280_loopback_sample_req_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_280_loopback_sample_req_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(20), ack => phi_stmt_280_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_entry_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(21) <= inputPort_3_Daemon_CP_407_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_entry_sample_req
      -- 
    phi_stmt_280_entry_sample_req_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_280_entry_sample_req_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(22), ack => phi_stmt_280_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_280_phi_mux_ack
      -- 
    phi_stmt_280_phi_mux_ack_452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_280_ack_0, ack => inputPort_3_Daemon_CP_407_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/type_cast_283_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/type_cast_283_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/type_cast_283_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/type_cast_283_sample_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/type_cast_283_update_start_
      -- CP-element group 25: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/type_cast_283_update_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/type_cast_283_update_completed__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(26) <= inputPort_3_Daemon_CP_407_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/type_cast_283_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(25), ack => inputPort_3_Daemon_CP_407_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_sample_start__ps
      -- 
    req_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(28), ack => next_count_down_317_284_buf_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_Update/req
      -- CP-element group 29: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_update_start_
      -- CP-element group 29: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_update_start__ps
      -- 
    req_478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(29), ack => next_count_down_317_284_buf_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_sample_completed__ps
      -- 
    ack_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_317_284_buf_ack_0, ack => inputPort_3_Daemon_CP_407_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_count_down_284_update_completed__ps
      -- 
    ack_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_317_284_buf_ack_1, ack => inputPort_3_Daemon_CP_407_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_285_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_sample_start_
      -- 
    rr_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(33), ack => RPIPE_in_data_3_287_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(11) & inputPort_3_Daemon_CP_407_elements(36);
      gj_inputPort_3_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_update_start_
      -- 
    cr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(34), ack => RPIPE_in_data_3_287_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(13) & inputPort_3_Daemon_CP_407_elements(35);
      gj_inputPort_3_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_sample_completed_
      -- 
    ra_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_3_287_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/RPIPE_in_data_3_287_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_285_update_completed_
      -- 
    ca_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_3_287_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_sample_start_
      -- 
    inputPort_3_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(12);
      gj_inputPort_3_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_sample_start__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(39) <= inputPort_3_Daemon_CP_407_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_sample_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_update_start__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(41) <= inputPort_3_Daemon_CP_407_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_update_completed__ps
      -- CP-element group 42: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_loopback_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(43) <= inputPort_3_Daemon_CP_407_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_loopback_sample_req_ps
      -- CP-element group 44: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_loopback_sample_req
      -- 
    phi_stmt_288_loopback_sample_req_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_288_loopback_sample_req_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(44), ack => phi_stmt_288_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_entry_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(45) <= inputPort_3_Daemon_CP_407_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_entry_sample_req_ps
      -- CP-element group 46: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_entry_sample_req
      -- 
    phi_stmt_288_entry_sample_req_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_288_entry_sample_req_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(46), ack => phi_stmt_288_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_phi_mux_ack_ps
      -- CP-element group 47: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/phi_stmt_288_phi_mux_ack
      -- 
    phi_stmt_288_phi_mux_ack_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_288_ack_0, ack => inputPort_3_Daemon_CP_407_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/konst_290_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/konst_290_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/konst_290_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/konst_290_sample_start_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/konst_290_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/konst_290_update_start_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/konst_290_update_completed__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(50) <= inputPort_3_Daemon_CP_407_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/konst_290_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(49), ack => inputPort_3_Daemon_CP_407_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_sample_start__ps
      -- 
    req_535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(52), ack => next_last_dest_id_323_291_buf_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_update_start_
      -- CP-element group 53: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_Update/req
      -- CP-element group 53: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_Update/$entry
      -- 
    req_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(53), ack => next_last_dest_id_323_291_buf_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_sample_completed__ps
      -- 
    ack_536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_323_291_buf_ack_0, ack => inputPort_3_Daemon_CP_407_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/R_next_last_dest_id_291_Update/$exit
      -- 
    ack_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_323_291_buf_ack_1, ack => inputPort_3_Daemon_CP_407_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_Sample/$entry
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(56), ack => WPIPE_noblock_obuf_3_1_335_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(58);
      gj_inputPort_3_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_Update/req
      -- CP-element group 57: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_update_start_
      -- CP-element group 57: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_sample_completed_
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_1_335_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(57)); -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(57), ack => WPIPE_noblock_obuf_3_1_335_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_1_335_update_completed_
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_1_335_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_Sample/req
      -- CP-element group 59: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_Sample/$entry
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(59), ack => WPIPE_noblock_obuf_3_2_344_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(61);
      gj_inputPort_3_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_Update/req
      -- CP-element group 60: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_update_start_
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_2_344_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(60)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(60), ack => WPIPE_noblock_obuf_3_2_344_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_Update/ack
      -- CP-element group 61: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_2_344_update_completed_
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_2_344_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_sample_start_
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(62), ack => WPIPE_noblock_obuf_3_3_353_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(64);
      gj_inputPort_3_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_Update/req
      -- CP-element group 63: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_update_start_
      -- CP-element group 63: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_sample_completed_
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_3_353_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(63)); -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(63), ack => WPIPE_noblock_obuf_3_3_353_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_3_353_Update/$exit
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_3_353_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_Sample/$entry
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(65), ack => WPIPE_noblock_obuf_3_4_362_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(67);
      gj_inputPort_3_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_Update/req
      -- CP-element group 66: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_update_start_
      -- CP-element group 66: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_Sample/$exit
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_4_362_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(66)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(66), ack => WPIPE_noblock_obuf_3_4_362_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/WPIPE_noblock_obuf_3_4_362_update_completed_
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_4_362_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(9), ack => inputPort_3_Daemon_CP_407_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_277/do_while_stmt_278/do_while_stmt_278_loop_body/$exit
      -- 
    inputPort_3_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(12) & inputPort_3_Daemon_CP_407_elements(58) & inputPort_3_Daemon_CP_407_elements(61) & inputPort_3_Daemon_CP_407_elements(64) & inputPort_3_Daemon_CP_407_elements(67);
      gj_inputPort_3_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_277/do_while_stmt_278/loop_exit/ack
      -- CP-element group 70: 	 branch_block_stmt_277/do_while_stmt_278/loop_exit/$exit
      -- 
    ack_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_278_branch_ack_0, ack => inputPort_3_Daemon_CP_407_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_277/do_while_stmt_278/loop_taken/ack
      -- CP-element group 71: 	 branch_block_stmt_277/do_while_stmt_278/loop_taken/$exit
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_278_branch_ack_1, ack => inputPort_3_Daemon_CP_407_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_277/do_while_stmt_278/$exit
      -- 
    inputPort_3_Daemon_CP_407_elements(72) <= inputPort_3_Daemon_CP_407_elements(3);
    inputPort_3_Daemon_do_while_stmt_278_terminator_608: loop_terminator -- 
      generic map (name => " inputPort_3_Daemon_do_while_stmt_278_terminator_608", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_3_Daemon_CP_407_elements(6),loop_continue => inputPort_3_Daemon_CP_407_elements(71),loop_terminate => inputPort_3_Daemon_CP_407_elements(70),loop_back => inputPort_3_Daemon_CP_407_elements(4),loop_exit => inputPort_3_Daemon_CP_407_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_280_phi_seq_480_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_3_Daemon_CP_407_elements(21);
      inputPort_3_Daemon_CP_407_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_3_Daemon_CP_407_elements(24);
      inputPort_3_Daemon_CP_407_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_3_Daemon_CP_407_elements(26);
      inputPort_3_Daemon_CP_407_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_3_Daemon_CP_407_elements(19);
      inputPort_3_Daemon_CP_407_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_3_Daemon_CP_407_elements(30);
      inputPort_3_Daemon_CP_407_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_3_Daemon_CP_407_elements(31);
      inputPort_3_Daemon_CP_407_elements(20) <= phi_mux_reqs(1);
      phi_stmt_280_phi_seq_480 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_280_phi_seq_480") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_3_Daemon_CP_407_elements(11), 
          phi_sample_ack => inputPort_3_Daemon_CP_407_elements(17), 
          phi_update_req => inputPort_3_Daemon_CP_407_elements(13), 
          phi_update_ack => inputPort_3_Daemon_CP_407_elements(18), 
          phi_mux_ack => inputPort_3_Daemon_CP_407_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_288_phi_seq_542_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_3_Daemon_CP_407_elements(45);
      inputPort_3_Daemon_CP_407_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_3_Daemon_CP_407_elements(48);
      inputPort_3_Daemon_CP_407_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_3_Daemon_CP_407_elements(50);
      inputPort_3_Daemon_CP_407_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_3_Daemon_CP_407_elements(43);
      inputPort_3_Daemon_CP_407_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_3_Daemon_CP_407_elements(54);
      inputPort_3_Daemon_CP_407_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_3_Daemon_CP_407_elements(55);
      inputPort_3_Daemon_CP_407_elements(44) <= phi_mux_reqs(1);
      phi_stmt_288_phi_seq_542 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_288_phi_seq_542") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_3_Daemon_CP_407_elements(39), 
          phi_sample_ack => inputPort_3_Daemon_CP_407_elements(40), 
          phi_update_req => inputPort_3_Daemon_CP_407_elements(41), 
          phi_update_ack => inputPort_3_Daemon_CP_407_elements(42), 
          phi_mux_ack => inputPort_3_Daemon_CP_407_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_432_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_3_Daemon_CP_407_elements(7);
        preds(1)  <= inputPort_3_Daemon_CP_407_elements(8);
        entry_tmerge_432 : transition_merge -- 
          generic map(name => " entry_tmerge_432")
          port map (preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_3_287_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_325_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_312_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_315_wire : std_logic_vector(15 downto 0);
    signal count_down_280 : std_logic_vector(15 downto 0);
    signal data_to_outport_328 : std_logic_vector(32 downto 0);
    signal dest_id_303 : std_logic_vector(7 downto 0);
    signal input_word_285 : std_logic_vector(31 downto 0);
    signal konst_290_wire_constant : std_logic_vector(7 downto 0);
    signal konst_295_wire_constant : std_logic_vector(15 downto 0);
    signal konst_311_wire_constant : std_logic_vector(15 downto 0);
    signal konst_314_wire_constant : std_logic_vector(15 downto 0);
    signal konst_331_wire_constant : std_logic_vector(7 downto 0);
    signal konst_340_wire_constant : std_logic_vector(7 downto 0);
    signal konst_349_wire_constant : std_logic_vector(7 downto 0);
    signal konst_358_wire_constant : std_logic_vector(7 downto 0);
    signal konst_376_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_288 : std_logic_vector(7 downto 0);
    signal new_packet_297 : std_logic_vector(0 downto 0);
    signal next_count_down_317 : std_logic_vector(15 downto 0);
    signal next_count_down_317_284_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_323 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_323_291_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_307 : std_logic_vector(15 downto 0);
    signal send_to_1_333 : std_logic_vector(0 downto 0);
    signal send_to_2_342 : std_logic_vector(0 downto 0);
    signal send_to_3_351 : std_logic_vector(0 downto 0);
    signal send_to_4_360 : std_logic_vector(0 downto 0);
    signal type_cast_283_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_325_wire_constant <= "1";
    konst_290_wire_constant <= "00000000";
    konst_295_wire_constant <= "0000000000000000";
    konst_311_wire_constant <= "0000000000000001";
    konst_314_wire_constant <= "0000000000000001";
    konst_331_wire_constant <= "00000001";
    konst_340_wire_constant <= "00000010";
    konst_349_wire_constant <= "00000011";
    konst_358_wire_constant <= "00000100";
    konst_376_wire_constant <= "1";
    type_cast_283_wire_constant <= "0000000000000000";
    phi_stmt_280: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_283_wire_constant & next_count_down_317_284_buffered;
      req <= phi_stmt_280_req_0 & phi_stmt_280_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_280",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_280_ack_0,
          idata => idata,
          odata => count_down_280,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_280
    phi_stmt_288: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_290_wire_constant & next_last_dest_id_323_291_buffered;
      req <= phi_stmt_288_req_0 & phi_stmt_288_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_288",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_288_ack_0,
          idata => idata,
          odata => last_dest_id_288,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_288
    -- flow-through select operator MUX_316_inst
    next_count_down_317 <= SUB_u16_u16_312_wire when (new_packet_297(0) /=  '0') else SUB_u16_u16_315_wire;
    -- flow-through select operator MUX_322_inst
    next_last_dest_id_323 <= dest_id_303 when (new_packet_297(0) /=  '0') else last_dest_id_288;
    -- flow-through slice operator slice_302_inst
    dest_id_303 <= input_word_285(31 downto 24);
    -- flow-through slice operator slice_306_inst
    pkt_length_307 <= input_word_285(23 downto 8);
    next_count_down_317_284_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_317_284_buf_req_0;
      next_count_down_317_284_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_317_284_buf_req_1;
      next_count_down_317_284_buf_ack_1<= rack(0);
      next_count_down_317_284_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_317_284_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_317_284_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_323_291_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_323_291_buf_req_0;
      next_last_dest_id_323_291_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_323_291_buf_req_1;
      next_last_dest_id_323_291_buf_ack_1<= rack(0);
      next_last_dest_id_323_291_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_323_291_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_323,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_323_291_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_285
    process(RPIPE_in_data_3_287_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_3_287_wire(31 downto 0);
      input_word_285 <= tmp_var; -- 
    end process;
    do_while_stmt_278_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_376_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_278_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_278_branch_req_0,
          ack0 => do_while_stmt_278_branch_ack_0,
          ack1 => do_while_stmt_278_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_327_inst
    process(R_ONE_1_325_wire_constant, input_word_285) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_325_wire_constant, input_word_285, tmp_var);
      data_to_outport_328 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_296_inst
    process(count_down_280) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_280, konst_295_wire_constant, tmp_var);
      new_packet_297 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_332_inst
    process(next_last_dest_id_323) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_323, konst_331_wire_constant, tmp_var);
      send_to_1_333 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_341_inst
    process(next_last_dest_id_323) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_323, konst_340_wire_constant, tmp_var);
      send_to_2_342 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_350_inst
    process(next_last_dest_id_323) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_323, konst_349_wire_constant, tmp_var);
      send_to_3_351 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_359_inst
    process(next_last_dest_id_323) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_323, konst_358_wire_constant, tmp_var);
      send_to_4_360 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_312_inst
    process(pkt_length_307) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_307, konst_311_wire_constant, tmp_var);
      SUB_u16_u16_312_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_315_inst
    process(count_down_280) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_280, konst_314_wire_constant, tmp_var);
      SUB_u16_u16_315_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_3_287_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_3_287_inst_req_0;
      RPIPE_in_data_3_287_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_3_287_inst_req_1;
      RPIPE_in_data_3_287_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_3_287_wire <= data_out(31 downto 0);
      in_data_3_read_0_gI: SplitGuardInterface generic map(name => "in_data_3_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_3_read_0: InputPortRevised -- 
        generic map ( name => "in_data_3_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_3_pipe_read_req(0),
          oack => in_data_3_pipe_read_ack(0),
          odata => in_data_3_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_3_1_335_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_1_335_inst_req_0;
      WPIPE_noblock_obuf_3_1_335_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_1_335_inst_req_1;
      WPIPE_noblock_obuf_3_1_335_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_333(0);
      data_in <= data_to_outport_328;
      noblock_obuf_3_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_1_pipe_write_req(0),
          oack => noblock_obuf_3_1_pipe_write_ack(0),
          odata => noblock_obuf_3_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_3_2_344_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_2_344_inst_req_0;
      WPIPE_noblock_obuf_3_2_344_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_2_344_inst_req_1;
      WPIPE_noblock_obuf_3_2_344_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_342(0);
      data_in <= data_to_outport_328;
      noblock_obuf_3_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_2_pipe_write_req(0),
          oack => noblock_obuf_3_2_pipe_write_ack(0),
          odata => noblock_obuf_3_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_3_3_353_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_3_353_inst_req_0;
      WPIPE_noblock_obuf_3_3_353_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_3_353_inst_req_1;
      WPIPE_noblock_obuf_3_3_353_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_351(0);
      data_in <= data_to_outport_328;
      noblock_obuf_3_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_3_pipe_write_req(0),
          oack => noblock_obuf_3_3_pipe_write_ack(0),
          odata => noblock_obuf_3_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_3_4_362_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_4_362_inst_req_0;
      WPIPE_noblock_obuf_3_4_362_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_4_362_inst_req_1;
      WPIPE_noblock_obuf_3_4_362_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_360(0);
      data_in <= data_to_outport_328;
      noblock_obuf_3_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_4_pipe_write_req(0),
          oack => noblock_obuf_3_4_pipe_write_ack(0),
          odata => noblock_obuf_3_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_3_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_4_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_4_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_4_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_4_Daemon;
architecture inputPort_4_Daemon_arch of inputPort_4_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_4_Daemon_CP_609_start: Boolean;
  signal inputPort_4_Daemon_CP_609_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_381_branch_req_0 : boolean;
  signal phi_stmt_383_req_1 : boolean;
  signal phi_stmt_383_req_0 : boolean;
  signal phi_stmt_383_ack_0 : boolean;
  signal next_count_down_420_387_buf_req_0 : boolean;
  signal next_count_down_420_387_buf_ack_0 : boolean;
  signal next_count_down_420_387_buf_req_1 : boolean;
  signal next_count_down_420_387_buf_ack_1 : boolean;
  signal RPIPE_in_data_4_390_inst_req_0 : boolean;
  signal RPIPE_in_data_4_390_inst_ack_0 : boolean;
  signal RPIPE_in_data_4_390_inst_req_1 : boolean;
  signal RPIPE_in_data_4_390_inst_ack_1 : boolean;
  signal phi_stmt_391_req_1 : boolean;
  signal phi_stmt_391_req_0 : boolean;
  signal phi_stmt_391_ack_0 : boolean;
  signal next_last_dest_id_426_394_buf_req_0 : boolean;
  signal next_last_dest_id_426_394_buf_ack_0 : boolean;
  signal next_last_dest_id_426_394_buf_req_1 : boolean;
  signal next_last_dest_id_426_394_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_1_438_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_1_438_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_1_438_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_1_438_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_2_447_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_2_447_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_2_447_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_2_447_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_456_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_3_456_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_3_456_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_456_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_4_465_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_465_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_465_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_4_465_inst_ack_1 : boolean;
  signal do_while_stmt_381_branch_ack_0 : boolean;
  signal do_while_stmt_381_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_4_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_4_Daemon_CP_609_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_4_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_4_Daemon_CP_609: Block -- control-path 
    signal inputPort_4_Daemon_CP_609_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_4_Daemon_CP_609_elements(0) <= inputPort_4_Daemon_CP_609_start;
    inputPort_4_Daemon_CP_609_symbol <= inputPort_4_Daemon_CP_609_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_380/branch_block_stmt_380__entry__
      -- CP-element group 0: 	 branch_block_stmt_380/do_while_stmt_381__entry__
      -- CP-element group 0: 	 branch_block_stmt_380/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_380/$exit
      -- CP-element group 1: 	 branch_block_stmt_380/branch_block_stmt_380__exit__
      -- CP-element group 1: 	 branch_block_stmt_380/do_while_stmt_381__exit__
      -- CP-element group 1: 	 $exit
      -- 
    inputPort_4_Daemon_CP_609_elements(1) <= inputPort_4_Daemon_CP_609_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381__entry__
      -- CP-element group 2: 	 branch_block_stmt_380/do_while_stmt_381/$entry
      -- 
    inputPort_4_Daemon_CP_609_elements(2) <= inputPort_4_Daemon_CP_609_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381__exit__
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_380/do_while_stmt_381/loop_back
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	71 
    -- CP-element group 5: 	70 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_380/do_while_stmt_381/condition_done
      -- CP-element group 5: 	 branch_block_stmt_380/do_while_stmt_381/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_380/do_while_stmt_381/loop_taken/$entry
      -- 
    inputPort_4_Daemon_CP_609_elements(5) <= inputPort_4_Daemon_CP_609_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_380/do_while_stmt_381/loop_body_done
      -- 
    inputPort_4_Daemon_CP_609_elements(6) <= inputPort_4_Daemon_CP_609_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/back_edge_to_loop_body
      -- 
    inputPort_4_Daemon_CP_609_elements(7) <= inputPort_4_Daemon_CP_609_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/first_time_through_loop_body
      -- 
    inputPort_4_Daemon_CP_609_elements(8) <= inputPort_4_Daemon_CP_609_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	68 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_388_sample_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	68 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/condition_evaluated
      -- 
    condition_evaluated_633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(10), ack => do_while_stmt_381_branch_req_0); -- 
    inputPort_4_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(68) & inputPort_4_Daemon_CP_609_elements(14);
      gj_inputPort_4_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_sample_start__ps
      -- 
    inputPort_4_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(15) & inputPort_4_Daemon_CP_609_elements(37) & inputPort_4_Daemon_CP_609_elements(14);
      gj_inputPort_4_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_388_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_sample_completed_
      -- 
    inputPort_4_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(17) & inputPort_4_Daemon_CP_609_elements(35) & inputPort_4_Daemon_CP_609_elements(40);
      gj_inputPort_4_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/aggregated_phi_update_req
      -- 
    inputPort_4_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(16) & inputPort_4_Daemon_CP_609_elements(32) & inputPort_4_Daemon_CP_609_elements(38);
      gj_inputPort_4_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_4_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42);
      gj_inputPort_4_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_sample_start_
      -- 
    inputPort_4_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(57) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(66);
      gj_inputPort_4_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_sample_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_update_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_loopback_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(19) <= inputPort_4_Daemon_CP_609_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_loopback_sample_req_ps
      -- 
    phi_stmt_383_loopback_sample_req_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_383_loopback_sample_req_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(20), ack => phi_stmt_383_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_entry_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(21) <= inputPort_4_Daemon_CP_609_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_entry_sample_req_ps
      -- 
    phi_stmt_383_entry_sample_req_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_383_entry_sample_req_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(22), ack => phi_stmt_383_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_383_phi_mux_ack_ps
      -- 
    phi_stmt_383_phi_mux_ack_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_383_ack_0, ack => inputPort_4_Daemon_CP_609_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/type_cast_386_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/type_cast_386_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/type_cast_386_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/type_cast_386_sample_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/type_cast_386_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/type_cast_386_update_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/type_cast_386_update_completed__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(26) <= inputPort_4_Daemon_CP_609_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/type_cast_386_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(25), ack => inputPort_4_Daemon_CP_609_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_Sample/req
      -- 
    req_675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(28), ack => next_count_down_420_387_buf_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_update_start_
      -- CP-element group 29: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_Update/req
      -- 
    req_680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(29), ack => next_count_down_420_387_buf_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_Sample/ack
      -- 
    ack_676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_420_387_buf_ack_0, ack => inputPort_4_Daemon_CP_609_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_count_down_387_Update/ack
      -- 
    ack_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_420_387_buf_ack_1, ack => inputPort_4_Daemon_CP_609_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_388_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(57) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(66);
      gj_inputPort_4_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_Sample/rr
      -- 
    rr_694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(33), ack => RPIPE_in_data_4_390_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(11) & inputPort_4_Daemon_CP_609_elements(36);
      gj_inputPort_4_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_update_start_
      -- CP-element group 34: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_Update/cr
      -- 
    cr_699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(34), ack => RPIPE_in_data_4_390_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(13) & inputPort_4_Daemon_CP_609_elements(35);
      gj_inputPort_4_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_Sample/ra
      -- 
    ra_695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_4_390_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_388_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/RPIPE_in_data_4_390_Update/ca
      -- 
    ca_700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_4_390_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_sample_start_
      -- 
    inputPort_4_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(57) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(66);
      gj_inputPort_4_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_sample_start__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(39) <= inputPort_4_Daemon_CP_609_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_sample_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_update_start__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(41) <= inputPort_4_Daemon_CP_609_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	14 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_update_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_loopback_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(43) <= inputPort_4_Daemon_CP_609_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_loopback_sample_req_ps
      -- 
    phi_stmt_391_loopback_sample_req_710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_391_loopback_sample_req_710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(44), ack => phi_stmt_391_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_entry_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(45) <= inputPort_4_Daemon_CP_609_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_entry_sample_req_ps
      -- 
    phi_stmt_391_entry_sample_req_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_391_entry_sample_req_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(46), ack => phi_stmt_391_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/phi_stmt_391_phi_mux_ack_ps
      -- 
    phi_stmt_391_phi_mux_ack_716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_391_ack_0, ack => inputPort_4_Daemon_CP_609_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/konst_393_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/konst_393_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/konst_393_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/konst_393_sample_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/konst_393_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/konst_393_update_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/konst_393_update_completed__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(50) <= inputPort_4_Daemon_CP_609_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/konst_393_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(49), ack => inputPort_4_Daemon_CP_609_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_Sample/req
      -- 
    req_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(52), ack => next_last_dest_id_426_394_buf_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_update_start_
      -- CP-element group 53: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_Update/req
      -- 
    req_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(53), ack => next_last_dest_id_426_394_buf_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_Sample/ack
      -- 
    ack_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_426_394_buf_ack_0, ack => inputPort_4_Daemon_CP_609_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/R_next_last_dest_id_394_Update/ack
      -- 
    ack_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_426_394_buf_ack_1, ack => inputPort_4_Daemon_CP_609_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_Sample/req
      -- 
    req_752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(56), ack => WPIPE_noblock_obuf_4_1_438_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(58);
      gj_inputPort_4_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_update_start_
      -- CP-element group 57: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_Update/req
      -- 
    ack_753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_1_438_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(57)); -- 
    req_757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(57), ack => WPIPE_noblock_obuf_4_1_438_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_1_438_Update/ack
      -- 
    ack_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_1_438_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_Sample/req
      -- 
    req_766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(59), ack => WPIPE_noblock_obuf_4_2_447_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(61);
      gj_inputPort_4_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_update_start_
      -- CP-element group 60: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_Update/req
      -- 
    ack_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_2_447_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(60)); -- 
    req_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(60), ack => WPIPE_noblock_obuf_4_2_447_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_2_447_Update/ack
      -- 
    ack_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_2_447_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_Sample/req
      -- 
    req_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(62), ack => WPIPE_noblock_obuf_4_3_456_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(64);
      gj_inputPort_4_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_update_start_
      -- CP-element group 63: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_Update/req
      -- 
    ack_781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_3_456_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(63)); -- 
    req_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(63), ack => WPIPE_noblock_obuf_4_3_456_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_3_456_Update/ack
      -- 
    ack_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_3_456_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_Sample/req
      -- 
    req_794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(65), ack => WPIPE_noblock_obuf_4_4_465_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(67);
      gj_inputPort_4_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_update_start_
      -- CP-element group 66: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_Update/req
      -- 
    ack_795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_4_465_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(66)); -- 
    req_799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(66), ack => WPIPE_noblock_obuf_4_4_465_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/WPIPE_noblock_obuf_4_4_465_Update/ack
      -- 
    ack_800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_4_465_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(9), ack => inputPort_4_Daemon_CP_609_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	12 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_380/do_while_stmt_381/do_while_stmt_381_loop_body/$exit
      -- 
    inputPort_4_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(64) & inputPort_4_Daemon_CP_609_elements(58) & inputPort_4_Daemon_CP_609_elements(67) & inputPort_4_Daemon_CP_609_elements(61) & inputPort_4_Daemon_CP_609_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_380/do_while_stmt_381/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_380/do_while_stmt_381/loop_exit/ack
      -- 
    ack_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_381_branch_ack_0, ack => inputPort_4_Daemon_CP_609_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_380/do_while_stmt_381/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_380/do_while_stmt_381/loop_taken/ack
      -- 
    ack_809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_381_branch_ack_1, ack => inputPort_4_Daemon_CP_609_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_380/do_while_stmt_381/$exit
      -- 
    inputPort_4_Daemon_CP_609_elements(72) <= inputPort_4_Daemon_CP_609_elements(3);
    inputPort_4_Daemon_do_while_stmt_381_terminator_810: loop_terminator -- 
      generic map (name => " inputPort_4_Daemon_do_while_stmt_381_terminator_810", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_4_Daemon_CP_609_elements(6),loop_continue => inputPort_4_Daemon_CP_609_elements(71),loop_terminate => inputPort_4_Daemon_CP_609_elements(70),loop_back => inputPort_4_Daemon_CP_609_elements(4),loop_exit => inputPort_4_Daemon_CP_609_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_383_phi_seq_682_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_4_Daemon_CP_609_elements(21);
      inputPort_4_Daemon_CP_609_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_4_Daemon_CP_609_elements(24);
      inputPort_4_Daemon_CP_609_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_4_Daemon_CP_609_elements(26);
      inputPort_4_Daemon_CP_609_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_4_Daemon_CP_609_elements(19);
      inputPort_4_Daemon_CP_609_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_4_Daemon_CP_609_elements(30);
      inputPort_4_Daemon_CP_609_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_4_Daemon_CP_609_elements(31);
      inputPort_4_Daemon_CP_609_elements(20) <= phi_mux_reqs(1);
      phi_stmt_383_phi_seq_682 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_383_phi_seq_682") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_4_Daemon_CP_609_elements(11), 
          phi_sample_ack => inputPort_4_Daemon_CP_609_elements(17), 
          phi_update_req => inputPort_4_Daemon_CP_609_elements(13), 
          phi_update_ack => inputPort_4_Daemon_CP_609_elements(18), 
          phi_mux_ack => inputPort_4_Daemon_CP_609_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_391_phi_seq_744_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_4_Daemon_CP_609_elements(45);
      inputPort_4_Daemon_CP_609_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_4_Daemon_CP_609_elements(48);
      inputPort_4_Daemon_CP_609_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_4_Daemon_CP_609_elements(50);
      inputPort_4_Daemon_CP_609_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_4_Daemon_CP_609_elements(43);
      inputPort_4_Daemon_CP_609_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_4_Daemon_CP_609_elements(54);
      inputPort_4_Daemon_CP_609_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_4_Daemon_CP_609_elements(55);
      inputPort_4_Daemon_CP_609_elements(44) <= phi_mux_reqs(1);
      phi_stmt_391_phi_seq_744 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_391_phi_seq_744") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_4_Daemon_CP_609_elements(39), 
          phi_sample_ack => inputPort_4_Daemon_CP_609_elements(40), 
          phi_update_req => inputPort_4_Daemon_CP_609_elements(41), 
          phi_update_ack => inputPort_4_Daemon_CP_609_elements(42), 
          phi_mux_ack => inputPort_4_Daemon_CP_609_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_634_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_4_Daemon_CP_609_elements(7);
        preds(1)  <= inputPort_4_Daemon_CP_609_elements(8);
        entry_tmerge_634 : transition_merge -- 
          generic map(name => " entry_tmerge_634")
          port map (preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_4_390_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_428_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_415_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_418_wire : std_logic_vector(15 downto 0);
    signal count_down_383 : std_logic_vector(15 downto 0);
    signal data_to_outport_431 : std_logic_vector(32 downto 0);
    signal dest_id_406 : std_logic_vector(7 downto 0);
    signal input_word_388 : std_logic_vector(31 downto 0);
    signal konst_393_wire_constant : std_logic_vector(7 downto 0);
    signal konst_398_wire_constant : std_logic_vector(15 downto 0);
    signal konst_414_wire_constant : std_logic_vector(15 downto 0);
    signal konst_417_wire_constant : std_logic_vector(15 downto 0);
    signal konst_434_wire_constant : std_logic_vector(7 downto 0);
    signal konst_443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_452_wire_constant : std_logic_vector(7 downto 0);
    signal konst_461_wire_constant : std_logic_vector(7 downto 0);
    signal konst_479_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_391 : std_logic_vector(7 downto 0);
    signal new_packet_400 : std_logic_vector(0 downto 0);
    signal next_count_down_420 : std_logic_vector(15 downto 0);
    signal next_count_down_420_387_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_426 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_426_394_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_410 : std_logic_vector(15 downto 0);
    signal send_to_1_436 : std_logic_vector(0 downto 0);
    signal send_to_2_445 : std_logic_vector(0 downto 0);
    signal send_to_3_454 : std_logic_vector(0 downto 0);
    signal send_to_4_463 : std_logic_vector(0 downto 0);
    signal type_cast_386_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_428_wire_constant <= "1";
    konst_393_wire_constant <= "00000000";
    konst_398_wire_constant <= "0000000000000000";
    konst_414_wire_constant <= "0000000000000001";
    konst_417_wire_constant <= "0000000000000001";
    konst_434_wire_constant <= "00000001";
    konst_443_wire_constant <= "00000010";
    konst_452_wire_constant <= "00000011";
    konst_461_wire_constant <= "00000100";
    konst_479_wire_constant <= "1";
    type_cast_386_wire_constant <= "0000000000000000";
    phi_stmt_383: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_386_wire_constant & next_count_down_420_387_buffered;
      req <= phi_stmt_383_req_0 & phi_stmt_383_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_383",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_383_ack_0,
          idata => idata,
          odata => count_down_383,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_383
    phi_stmt_391: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_393_wire_constant & next_last_dest_id_426_394_buffered;
      req <= phi_stmt_391_req_0 & phi_stmt_391_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_391",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_391_ack_0,
          idata => idata,
          odata => last_dest_id_391,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_391
    -- flow-through select operator MUX_419_inst
    next_count_down_420 <= SUB_u16_u16_415_wire when (new_packet_400(0) /=  '0') else SUB_u16_u16_418_wire;
    -- flow-through select operator MUX_425_inst
    next_last_dest_id_426 <= dest_id_406 when (new_packet_400(0) /=  '0') else last_dest_id_391;
    -- flow-through slice operator slice_405_inst
    dest_id_406 <= input_word_388(31 downto 24);
    -- flow-through slice operator slice_409_inst
    pkt_length_410 <= input_word_388(23 downto 8);
    next_count_down_420_387_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_420_387_buf_req_0;
      next_count_down_420_387_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_420_387_buf_req_1;
      next_count_down_420_387_buf_ack_1<= rack(0);
      next_count_down_420_387_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_420_387_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_420_387_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_426_394_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_426_394_buf_req_0;
      next_last_dest_id_426_394_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_426_394_buf_req_1;
      next_last_dest_id_426_394_buf_ack_1<= rack(0);
      next_last_dest_id_426_394_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_426_394_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_426,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_426_394_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_388
    process(RPIPE_in_data_4_390_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_4_390_wire(31 downto 0);
      input_word_388 <= tmp_var; -- 
    end process;
    do_while_stmt_381_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_479_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_381_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_381_branch_req_0,
          ack0 => do_while_stmt_381_branch_ack_0,
          ack1 => do_while_stmt_381_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_430_inst
    process(R_ONE_1_428_wire_constant, input_word_388) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_428_wire_constant, input_word_388, tmp_var);
      data_to_outport_431 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_399_inst
    process(count_down_383) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_383, konst_398_wire_constant, tmp_var);
      new_packet_400 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_435_inst
    process(next_last_dest_id_426) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_426, konst_434_wire_constant, tmp_var);
      send_to_1_436 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_444_inst
    process(next_last_dest_id_426) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_426, konst_443_wire_constant, tmp_var);
      send_to_2_445 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_453_inst
    process(next_last_dest_id_426) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_426, konst_452_wire_constant, tmp_var);
      send_to_3_454 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_462_inst
    process(next_last_dest_id_426) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_426, konst_461_wire_constant, tmp_var);
      send_to_4_463 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_415_inst
    process(pkt_length_410) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_410, konst_414_wire_constant, tmp_var);
      SUB_u16_u16_415_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_418_inst
    process(count_down_383) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_383, konst_417_wire_constant, tmp_var);
      SUB_u16_u16_418_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_4_390_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_4_390_inst_req_0;
      RPIPE_in_data_4_390_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_4_390_inst_req_1;
      RPIPE_in_data_4_390_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_4_390_wire <= data_out(31 downto 0);
      in_data_4_read_0_gI: SplitGuardInterface generic map(name => "in_data_4_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_4_read_0: InputPortRevised -- 
        generic map ( name => "in_data_4_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_4_pipe_read_req(0),
          oack => in_data_4_pipe_read_ack(0),
          odata => in_data_4_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_4_1_438_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_1_438_inst_req_0;
      WPIPE_noblock_obuf_4_1_438_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_1_438_inst_req_1;
      WPIPE_noblock_obuf_4_1_438_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_436(0);
      data_in <= data_to_outport_431;
      noblock_obuf_4_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_1_pipe_write_req(0),
          oack => noblock_obuf_4_1_pipe_write_ack(0),
          odata => noblock_obuf_4_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_4_2_447_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_2_447_inst_req_0;
      WPIPE_noblock_obuf_4_2_447_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_2_447_inst_req_1;
      WPIPE_noblock_obuf_4_2_447_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_445(0);
      data_in <= data_to_outport_431;
      noblock_obuf_4_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_2_pipe_write_req(0),
          oack => noblock_obuf_4_2_pipe_write_ack(0),
          odata => noblock_obuf_4_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_4_3_456_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_3_456_inst_req_0;
      WPIPE_noblock_obuf_4_3_456_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_3_456_inst_req_1;
      WPIPE_noblock_obuf_4_3_456_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_454(0);
      data_in <= data_to_outport_431;
      noblock_obuf_4_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_3_pipe_write_req(0),
          oack => noblock_obuf_4_3_pipe_write_ack(0),
          odata => noblock_obuf_4_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_4_4_465_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_4_465_inst_req_0;
      WPIPE_noblock_obuf_4_4_465_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_4_465_inst_req_1;
      WPIPE_noblock_obuf_4_4_465_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_463(0);
      data_in <= data_to_outport_431;
      noblock_obuf_4_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_4_pipe_write_req(0),
          oack => noblock_obuf_4_4_pipe_write_ack(0),
          odata => noblock_obuf_4_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_4_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_1_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_1_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_1_Daemon;
architecture outputPort_1_Daemon_arch of outputPort_1_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_1_Daemon_CP_814_start: Boolean;
  signal outputPort_1_Daemon_CP_814_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(15 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_with_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_with_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal RPIPE_noblock_obuf_2_1_670_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_1_1_665_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_670_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_665_inst_ack_1 : boolean;
  signal phi_stmt_661_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_670_inst_req_1 : boolean;
  signal phi_stmt_671_req_0 : boolean;
  signal phi_stmt_671_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_670_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_665_inst_req_0 : boolean;
  signal phi_stmt_666_req_1 : boolean;
  signal phi_stmt_661_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_665_inst_req_1 : boolean;
  signal phi_stmt_671_req_1 : boolean;
  signal phi_stmt_661_req_1 : boolean;
  signal phi_stmt_666_ack_0 : boolean;
  signal phi_stmt_666_req_0 : boolean;
  signal do_while_stmt_659_branch_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_675_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_675_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_675_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_1_675_inst_ack_1 : boolean;
  signal phi_stmt_676_req_1 : boolean;
  signal phi_stmt_676_req_0 : boolean;
  signal phi_stmt_676_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_680_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_680_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_680_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_1_680_inst_ack_1 : boolean;
  signal phi_stmt_681_req_1 : boolean;
  signal phi_stmt_681_req_0 : boolean;
  signal phi_stmt_681_ack_0 : boolean;
  signal next_active_packet_764_684_buf_req_0 : boolean;
  signal next_active_packet_764_684_buf_ack_0 : boolean;
  signal next_active_packet_764_684_buf_req_1 : boolean;
  signal next_active_packet_764_684_buf_ack_1 : boolean;
  signal phi_stmt_685_req_1 : boolean;
  signal phi_stmt_685_req_0 : boolean;
  signal phi_stmt_685_ack_0 : boolean;
  signal next_down_counter_819_688_buf_req_0 : boolean;
  signal next_down_counter_819_688_buf_ack_0 : boolean;
  signal next_down_counter_819_688_buf_req_1 : boolean;
  signal next_down_counter_819_688_buf_ack_1 : boolean;
  signal phi_stmt_689_req_1 : boolean;
  signal phi_stmt_689_req_0 : boolean;
  signal phi_stmt_689_ack_0 : boolean;
  signal next_pkt_with_priority_764_692_buf_req_0 : boolean;
  signal next_pkt_with_priority_764_692_buf_ack_0 : boolean;
  signal next_pkt_with_priority_764_692_buf_req_1 : boolean;
  signal next_pkt_with_priority_764_692_buf_ack_1 : boolean;
  signal WPIPE_out_data_1_904_inst_req_0 : boolean;
  signal WPIPE_out_data_1_904_inst_ack_0 : boolean;
  signal WPIPE_out_data_1_904_inst_req_1 : boolean;
  signal WPIPE_out_data_1_904_inst_ack_1 : boolean;
  signal do_while_stmt_659_branch_ack_0 : boolean;
  signal do_while_stmt_659_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_1_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_1_Daemon_CP_814_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_1_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_1_Daemon_CP_814: Block -- control-path 
    signal outputPort_1_Daemon_CP_814_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_1_Daemon_CP_814_elements(0) <= outputPort_1_Daemon_CP_814_start;
    outputPort_1_Daemon_CP_814_symbol <= outputPort_1_Daemon_CP_814_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_658/branch_block_stmt_658__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_658/$entry
      -- CP-element group 0: 	 branch_block_stmt_658/do_while_stmt_659__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_658/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_658/branch_block_stmt_658__exit__
      -- CP-element group 1: 	 branch_block_stmt_658/do_while_stmt_659__exit__
      -- 
    outputPort_1_Daemon_CP_814_elements(1) <= outputPort_1_Daemon_CP_814_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659__entry__
      -- CP-element group 2: 	 branch_block_stmt_658/do_while_stmt_659/$entry
      -- 
    outputPort_1_Daemon_CP_814_elements(2) <= outputPort_1_Daemon_CP_814_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659__exit__
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_658/do_while_stmt_659/loop_back
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	160 
    -- CP-element group 5: 	159 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_658/do_while_stmt_659/condition_done
      -- CP-element group 5: 	 branch_block_stmt_658/do_while_stmt_659/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_658/do_while_stmt_659/loop_taken/$entry
      -- 
    outputPort_1_Daemon_CP_814_elements(5) <= outputPort_1_Daemon_CP_814_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_658/do_while_stmt_659/loop_body_done
      -- 
    outputPort_1_Daemon_CP_814_elements(6) <= outputPort_1_Daemon_CP_814_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	104 
    -- CP-element group 7: 	122 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	42 
    -- CP-element group 7: 	63 
    -- CP-element group 7: 	84 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/back_edge_to_loop_body
      -- 
    outputPort_1_Daemon_CP_814_elements(7) <= outputPort_1_Daemon_CP_814_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	106 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	124 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	44 
    -- CP-element group 8: 	65 
    -- CP-element group 8: 	86 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/first_time_through_loop_body
      -- 
    outputPort_1_Daemon_CP_814_elements(8) <= outputPort_1_Daemon_CP_814_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	135 
    -- CP-element group 9: 	117 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	57 
    -- CP-element group 9: 	58 
    -- CP-element group 9: 	78 
    -- CP-element group 9: 	79 
    -- CP-element group 9: 	99 
    -- CP-element group 9: 	100 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/loop_body_start
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/condition_evaluated
      -- 
    condition_evaluated_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(10), ack => do_while_stmt_659_branch_req_0); -- 
    outputPort_1_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(157) & outputPort_1_Daemon_CP_814_elements(14);
      gj_outputPort_1_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	135 
    -- CP-element group 11: 	117 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11: 	99 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	101 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	38 
    -- CP-element group 11: 	59 
    -- CP-element group 11: 	80 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_sample_start__ps
      -- 
    outputPort_1_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(135) & outputPort_1_Daemon_CP_814_elements(117) & outputPort_1_Daemon_CP_814_elements(15) & outputPort_1_Daemon_CP_814_elements(36) & outputPort_1_Daemon_CP_814_elements(57) & outputPort_1_Daemon_CP_814_elements(78) & outputPort_1_Daemon_CP_814_elements(99) & outputPort_1_Daemon_CP_814_elements(14);
      gj_outputPort_1_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	102 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	138 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	39 
    -- CP-element group 12: 	60 
    -- CP-element group 12: 	81 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	135 
    -- CP-element group 12: 	117 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	57 
    -- CP-element group 12: 	78 
    -- CP-element group 12: 	99 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_sample_completed_
      -- 
    outputPort_1_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(102) & outputPort_1_Daemon_CP_814_elements(119) & outputPort_1_Daemon_CP_814_elements(138) & outputPort_1_Daemon_CP_814_elements(18) & outputPort_1_Daemon_CP_814_elements(39) & outputPort_1_Daemon_CP_814_elements(60) & outputPort_1_Daemon_CP_814_elements(81);
      gj_outputPort_1_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	136 
    -- CP-element group 13: 	118 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	58 
    -- CP-element group 13: 	79 
    -- CP-element group 13: 	100 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	139 
    -- CP-element group 13: 	120 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	40 
    -- CP-element group 13: 	61 
    -- CP-element group 13: 	82 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_update_start__ps
      -- 
    outputPort_1_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(136) & outputPort_1_Daemon_CP_814_elements(118) & outputPort_1_Daemon_CP_814_elements(16) & outputPort_1_Daemon_CP_814_elements(37) & outputPort_1_Daemon_CP_814_elements(58) & outputPort_1_Daemon_CP_814_elements(79) & outputPort_1_Daemon_CP_814_elements(100);
      gj_outputPort_1_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	103 
    -- CP-element group 14: 	121 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	41 
    -- CP-element group 14: 	62 
    -- CP-element group 14: 	83 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_1_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(140) & outputPort_1_Daemon_CP_814_elements(103) & outputPort_1_Daemon_CP_814_elements(121) & outputPort_1_Daemon_CP_814_elements(20) & outputPort_1_Daemon_CP_814_elements(41) & outputPort_1_Daemon_CP_814_elements(62) & outputPort_1_Daemon_CP_814_elements(83);
      gj_outputPort_1_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(17) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(19) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(21) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_loopback_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_loopback_sample_req
      -- 
    phi_stmt_661_loopback_sample_req_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_661_loopback_sample_req_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(22), ack => phi_stmt_661_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(23) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_entry_sample_req_ps
      -- CP-element group 24: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_entry_sample_req
      -- 
    phi_stmt_661_entry_sample_req_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_661_entry_sample_req_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(24), ack => phi_stmt_661_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_661_phi_mux_ack_ps
      -- 
    phi_stmt_661_phi_mux_ack_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_661_ack_0, ack => outputPort_1_Daemon_CP_814_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_663_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_663_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_663_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_663_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_663_update_start_
      -- CP-element group 27: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_663_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_663_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(28) <= outputPort_1_Daemon_CP_814_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_663_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(27), ack => outputPort_1_Daemon_CP_814_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	35 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_sample_start_
      -- 
    rr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(32), ack => RPIPE_noblock_obuf_1_1_665_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(30) & outputPort_1_Daemon_CP_814_elements(35);
      gj_outputPort_1_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: 	34 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_update_start_
      -- CP-element group 33: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_Update/cr
      -- 
    cr_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(33), ack => RPIPE_noblock_obuf_1_1_665_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(31) & outputPort_1_Daemon_CP_814_elements(34);
      gj_outputPort_1_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	33 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_sample_completed__ps
      -- 
    ra_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_1_665_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	32 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_1_1_665_update_completed__ps
      -- 
    ca_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_1_665_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	11 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	155 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	11 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(38) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	12 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	13 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(40) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	154 
    -- CP-element group 41: 	14 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	7 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(42) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_loopback_sample_req_ps
      -- 
    phi_stmt_666_loopback_sample_req_897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_666_loopback_sample_req_897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(43), ack => phi_stmt_666_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	8 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(44) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_entry_sample_req_ps
      -- CP-element group 45: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_entry_sample_req
      -- 
    phi_stmt_666_entry_sample_req_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_666_entry_sample_req_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(45), ack => phi_stmt_666_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_phi_mux_ack_ps
      -- CP-element group 46: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_666_phi_mux_ack
      -- 
    phi_stmt_666_phi_mux_ack_903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_666_ack_0, ack => outputPort_1_Daemon_CP_814_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_668_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_668_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_668_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_668_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_668_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_668_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_668_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(49) <= outputPort_1_Daemon_CP_814_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_668_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(48), ack => outputPort_1_Daemon_CP_814_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_Sample/$entry
      -- 
    rr_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(53), ack => RPIPE_noblock_obuf_2_1_670_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(51) & outputPort_1_Daemon_CP_814_elements(56);
      gj_outputPort_1_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: 	55 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_Update/cr
      -- CP-element group 54: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_update_start_
      -- 
    cr_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(54), ack => RPIPE_noblock_obuf_2_1_670_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(52) & outputPort_1_Daemon_CP_814_elements(55);
      gj_outputPort_1_Daemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	54 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_Sample/$exit
      -- 
    ra_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_1_670_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_2_1_670_update_completed_
      -- 
    ca_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_1_670_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(56)); -- 
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	9 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	12 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	11 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	9 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	155 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	13 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	11 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(59) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	12 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	13 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(61) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	154 
    -- CP-element group 62: 	14 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	7 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(63) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_loopback_sample_req_ps
      -- CP-element group 64: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_loopback_sample_req
      -- 
    phi_stmt_671_loopback_sample_req_941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_671_loopback_sample_req_941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(64), ack => phi_stmt_671_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	8 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(65) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_entry_sample_req_ps
      -- CP-element group 66: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_entry_sample_req
      -- 
    phi_stmt_671_entry_sample_req_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_671_entry_sample_req_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(66), ack => phi_stmt_671_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_phi_mux_ack
      -- CP-element group 67: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_671_phi_mux_ack_ps
      -- 
    phi_stmt_671_phi_mux_ack_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_671_ack_0, ack => outputPort_1_Daemon_CP_814_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_673_sample_start__ps
      -- CP-element group 68: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_673_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_673_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_673_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_673_update_start__ps
      -- CP-element group 69: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_673_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_673_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(70) <= outputPort_1_Daemon_CP_814_elements(71);
    -- CP-element group 71:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	70 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_673_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(69), ack => outputPort_1_Daemon_CP_814_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	77 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_Sample/rr
      -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(74), ack => RPIPE_noblock_obuf_3_1_675_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(72) & outputPort_1_Daemon_CP_814_elements(77);
      gj_outputPort_1_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	76 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_update_start_
      -- CP-element group 75: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_Update/cr
      -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(75), ack => RPIPE_noblock_obuf_3_1_675_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(73) & outputPort_1_Daemon_CP_814_elements(76);
      gj_outputPort_1_Daemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	75 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_Sample/ra
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_1_675_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(76)); -- 
    -- CP-element group 77:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	74 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_3_1_675_Update/ca
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_1_675_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	12 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	11 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	9 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	155 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	13 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	11 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(80) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 81:  join  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	12 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	13 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(82) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	154 
    -- CP-element group 83: 	14 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	7 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(84) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_loopback_sample_req
      -- CP-element group 85: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_loopback_sample_req_ps
      -- 
    phi_stmt_676_loopback_sample_req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_loopback_sample_req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(85), ack => phi_stmt_676_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	8 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(86) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 87:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_entry_sample_req
      -- CP-element group 87: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_entry_sample_req_ps
      -- 
    phi_stmt_676_entry_sample_req_988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_entry_sample_req_988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(87), ack => phi_stmt_676_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_phi_mux_ack
      -- CP-element group 88: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_676_phi_mux_ack_ps
      -- 
    phi_stmt_676_phi_mux_ack_991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_676_ack_0, ack => outputPort_1_Daemon_CP_814_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_678_sample_start__ps
      -- CP-element group 89: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_678_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_678_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_678_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_678_update_start__ps
      -- CP-element group 90: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_678_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_678_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(91) <= outputPort_1_Daemon_CP_814_elements(92);
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_33_678_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(90), ack => outputPort_1_Daemon_CP_814_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	98 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_Sample/rr
      -- 
    rr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(95), ack => RPIPE_noblock_obuf_4_1_680_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(93) & outputPort_1_Daemon_CP_814_elements(98);
      gj_outputPort_1_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	97 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_update_start_
      -- CP-element group 96: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_Update/cr
      -- 
    cr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(96), ack => RPIPE_noblock_obuf_4_1_680_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(94) & outputPort_1_Daemon_CP_814_elements(97);
      gj_outputPort_1_Daemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	96 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_sample_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_Sample/ra
      -- 
    ra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_1_680_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(97)); -- 
    -- CP-element group 98:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	95 
    -- CP-element group 98:  members (4) 
      -- CP-element group 98: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_update_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/RPIPE_noblock_obuf_4_1_680_Update/ca
      -- 
    ca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_1_680_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(98)); -- 
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	9 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	12 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	11 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	9 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	155 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	13 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	11 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(101) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	12 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	154 
    -- CP-element group 103: 	14 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(103) is bound as output of CP function.
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	7 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(104) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 105:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_loopback_sample_req
      -- CP-element group 105: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_loopback_sample_req_ps
      -- 
    phi_stmt_681_loopback_sample_req_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_loopback_sample_req_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(105), ack => phi_stmt_681_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	8 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(106) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 107:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_entry_sample_req
      -- CP-element group 107: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_entry_sample_req_ps
      -- 
    phi_stmt_681_entry_sample_req_1032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_entry_sample_req_1032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(107), ack => phi_stmt_681_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_phi_mux_ack
      -- CP-element group 108: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_681_phi_mux_ack_ps
      -- 
    phi_stmt_681_phi_mux_ack_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_681_ack_0, ack => outputPort_1_Daemon_CP_814_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_3_683_sample_start__ps
      -- CP-element group 109: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_3_683_sample_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_3_683_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_3_683_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_3_683_update_start__ps
      -- CP-element group 110: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_3_683_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_3_683_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(111) <= outputPort_1_Daemon_CP_814_elements(112);
    -- CP-element group 112:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	111 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_3_683_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(110), ack => outputPort_1_Daemon_CP_814_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_sample_start__ps
      -- CP-element group 113: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_Sample/req
      -- 
    req_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(113), ack => next_active_packet_764_684_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_update_start__ps
      -- CP-element group 114: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_update_start_
      -- CP-element group 114: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_Update/req
      -- 
    req_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(114), ack => next_active_packet_764_684_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_sample_completed__ps
      -- CP-element group 115: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_Sample/ack
      -- 
    ack_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_764_684_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(115)); -- 
    -- CP-element group 116:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_update_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_active_packet_684_Update/ack
      -- 
    ack_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_764_684_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(116)); -- 
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	9 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	12 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	11 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	155 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	13 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	12 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	13 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(120) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	154 
    -- CP-element group 121: 	14 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	7 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(122) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_loopback_sample_req
      -- CP-element group 123: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_loopback_sample_req_ps
      -- 
    phi_stmt_685_loopback_sample_req_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_685_loopback_sample_req_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(123), ack => phi_stmt_685_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(124) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_entry_sample_req
      -- CP-element group 125: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_entry_sample_req_ps
      -- 
    phi_stmt_685_entry_sample_req_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_685_entry_sample_req_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(125), ack => phi_stmt_685_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_phi_mux_ack
      -- CP-element group 126: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_685_phi_mux_ack_ps
      -- 
    phi_stmt_685_phi_mux_ack_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_685_ack_0, ack => outputPort_1_Daemon_CP_814_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_16_687_sample_start__ps
      -- CP-element group 127: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_16_687_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_16_687_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_16_687_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_16_687_update_start__ps
      -- CP-element group 128: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_16_687_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_16_687_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(129) <= outputPort_1_Daemon_CP_814_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_ZERO_16_687_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(128), ack => outputPort_1_Daemon_CP_814_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_sample_start__ps
      -- CP-element group 131: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_Sample/req
      -- 
    req_1100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(131), ack => next_down_counter_819_688_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_update_start__ps
      -- CP-element group 132: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_update_start_
      -- CP-element group 132: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_Update/req
      -- 
    req_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(132), ack => next_down_counter_819_688_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_Sample/ack
      -- 
    ack_1101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_819_688_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(133)); -- 
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_down_counter_688_Update/ack
      -- 
    ack_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_819_688_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	9 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	11 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	155 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	13 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(137) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	12 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	13 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(139) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(141) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_loopback_sample_req_ps
      -- 
    phi_stmt_689_loopback_sample_req_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_689_loopback_sample_req_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(142), ack => phi_stmt_689_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(143) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_entry_sample_req_ps
      -- 
    phi_stmt_689_entry_sample_req_1120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_689_entry_sample_req_1120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(144), ack => phi_stmt_689_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/phi_stmt_689_phi_mux_ack_ps
      -- 
    phi_stmt_689_phi_mux_ack_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_689_ack_0, ack => outputPort_1_Daemon_CP_814_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/konst_691_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/konst_691_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/konst_691_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/konst_691_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/konst_691_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/konst_691_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/konst_691_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(148) <= outputPort_1_Daemon_CP_814_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/konst_691_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(147), ack => outputPort_1_Daemon_CP_814_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_Sample/req
      -- 
    req_1144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(150), ack => next_pkt_with_priority_764_692_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_update_start_
      -- CP-element group 151: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_Update/req
      -- 
    req_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(151), ack => next_pkt_with_priority_764_692_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_Sample/ack
      -- 
    ack_1145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_with_priority_764_692_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/R_next_pkt_with_priority_692_Update/ack
      -- 
    ack_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_with_priority_764_692_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	103 
    -- CP-element group 154: 	121 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	41 
    -- CP-element group 154: 	62 
    -- CP-element group 154: 	83 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_Sample/req
      -- 
    req_1159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(154), ack => WPIPE_out_data_1_904_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(140) & outputPort_1_Daemon_CP_814_elements(103) & outputPort_1_Daemon_CP_814_elements(121) & outputPort_1_Daemon_CP_814_elements(20) & outputPort_1_Daemon_CP_814_elements(41) & outputPort_1_Daemon_CP_814_elements(62) & outputPort_1_Daemon_CP_814_elements(83) & outputPort_1_Daemon_CP_814_elements(156);
      gj_outputPort_1_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	136 
    -- CP-element group 155: 	118 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	37 
    -- CP-element group 155: 	58 
    -- CP-element group 155: 	79 
    -- CP-element group 155: 	100 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_update_start_
      -- CP-element group 155: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_Update/req
      -- 
    ack_1160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_1_904_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(155)); -- 
    req_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(155), ack => WPIPE_out_data_1_904_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/WPIPE_out_data_1_904_Update/ack
      -- 
    ack_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_1_904_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(9), ack => outputPort_1_Daemon_CP_814_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_658/do_while_stmt_659/do_while_stmt_659_loop_body/$exit
      -- 
    outputPort_1_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(156) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_658/do_while_stmt_659/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_658/do_while_stmt_659/loop_exit/ack
      -- 
    ack_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_659_branch_ack_0, ack => outputPort_1_Daemon_CP_814_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_658/do_while_stmt_659/loop_taken/$exit
      -- CP-element group 160: 	 branch_block_stmt_658/do_while_stmt_659/loop_taken/ack
      -- 
    ack_1174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_659_branch_ack_1, ack => outputPort_1_Daemon_CP_814_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_658/do_while_stmt_659/$exit
      -- 
    outputPort_1_Daemon_CP_814_elements(161) <= outputPort_1_Daemon_CP_814_elements(3);
    outputPort_1_Daemon_do_while_stmt_659_terminator_1175: loop_terminator -- 
      generic map (name => " outputPort_1_Daemon_do_while_stmt_659_terminator_1175", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_1_Daemon_CP_814_elements(6),loop_continue => outputPort_1_Daemon_CP_814_elements(160),loop_terminate => outputPort_1_Daemon_CP_814_elements(159),loop_back => outputPort_1_Daemon_CP_814_elements(4),loop_exit => outputPort_1_Daemon_CP_814_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_661_phi_seq_887_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(23);
      outputPort_1_Daemon_CP_814_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(26);
      outputPort_1_Daemon_CP_814_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(28);
      outputPort_1_Daemon_CP_814_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(21);
      outputPort_1_Daemon_CP_814_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(34);
      outputPort_1_Daemon_CP_814_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(35);
      outputPort_1_Daemon_CP_814_elements(22) <= phi_mux_reqs(1);
      phi_stmt_661_phi_seq_887 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_661_phi_seq_887") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(17), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(18), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(19), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(20), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_666_phi_seq_931_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(44);
      outputPort_1_Daemon_CP_814_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(47);
      outputPort_1_Daemon_CP_814_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(49);
      outputPort_1_Daemon_CP_814_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(42);
      outputPort_1_Daemon_CP_814_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(55);
      outputPort_1_Daemon_CP_814_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(56);
      outputPort_1_Daemon_CP_814_elements(43) <= phi_mux_reqs(1);
      phi_stmt_666_phi_seq_931 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_666_phi_seq_931") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(38), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(39), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(40), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(41), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_671_phi_seq_975_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(65);
      outputPort_1_Daemon_CP_814_elements(68)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(68);
      outputPort_1_Daemon_CP_814_elements(69)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(70);
      outputPort_1_Daemon_CP_814_elements(66) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(63);
      outputPort_1_Daemon_CP_814_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(76);
      outputPort_1_Daemon_CP_814_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(77);
      outputPort_1_Daemon_CP_814_elements(64) <= phi_mux_reqs(1);
      phi_stmt_671_phi_seq_975 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_671_phi_seq_975") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(59), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(60), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(61), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(62), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(67), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_676_phi_seq_1019_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(86);
      outputPort_1_Daemon_CP_814_elements(89)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(89);
      outputPort_1_Daemon_CP_814_elements(90)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(91);
      outputPort_1_Daemon_CP_814_elements(87) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(84);
      outputPort_1_Daemon_CP_814_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(97);
      outputPort_1_Daemon_CP_814_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(98);
      outputPort_1_Daemon_CP_814_elements(85) <= phi_mux_reqs(1);
      phi_stmt_676_phi_seq_1019 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_676_phi_seq_1019") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(80), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(81), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(82), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(83), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(88), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_681_phi_seq_1063_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(106);
      outputPort_1_Daemon_CP_814_elements(109)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(109);
      outputPort_1_Daemon_CP_814_elements(110)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(111);
      outputPort_1_Daemon_CP_814_elements(107) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(104);
      outputPort_1_Daemon_CP_814_elements(113)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(115);
      outputPort_1_Daemon_CP_814_elements(114)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(116);
      outputPort_1_Daemon_CP_814_elements(105) <= phi_mux_reqs(1);
      phi_stmt_681_phi_seq_1063 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_681_phi_seq_1063") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(101), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(102), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(13), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(103), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(108), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_685_phi_seq_1107_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(124);
      outputPort_1_Daemon_CP_814_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(127);
      outputPort_1_Daemon_CP_814_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(129);
      outputPort_1_Daemon_CP_814_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(122);
      outputPort_1_Daemon_CP_814_elements(131)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(133);
      outputPort_1_Daemon_CP_814_elements(132)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(134);
      outputPort_1_Daemon_CP_814_elements(123) <= phi_mux_reqs(1);
      phi_stmt_685_phi_seq_1107 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_685_phi_seq_1107") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(11), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(119), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(120), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(121), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_689_phi_seq_1151_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(143);
      outputPort_1_Daemon_CP_814_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(146);
      outputPort_1_Daemon_CP_814_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(148);
      outputPort_1_Daemon_CP_814_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(141);
      outputPort_1_Daemon_CP_814_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(152);
      outputPort_1_Daemon_CP_814_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(153);
      outputPort_1_Daemon_CP_814_elements(142) <= phi_mux_reqs(1);
      phi_stmt_689_phi_seq_1151 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_689_phi_seq_1151") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(137), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(138), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(139), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(140), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_839_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_1_Daemon_CP_814_elements(7);
        preds(1)  <= outputPort_1_Daemon_CP_814_elements(8);
        entry_tmerge_839 : transition_merge -- 
          generic map(name => " entry_tmerge_839")
          port map (preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u16_u1_804_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_729_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_735_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_742_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_748_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_768_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_775_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_783_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_790_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_825_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_833_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_841_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_849_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_855_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_860_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_865_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_877_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_883_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_890_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_896_wire : std_logic_vector(0 downto 0);
    signal MUX_732_wire : std_logic_vector(0 downto 0);
    signal MUX_738_wire : std_logic_vector(0 downto 0);
    signal MUX_745_wire : std_logic_vector(0 downto 0);
    signal MUX_751_wire : std_logic_vector(0 downto 0);
    signal MUX_772_wire : std_logic_vector(15 downto 0);
    signal MUX_779_wire : std_logic_vector(15 downto 0);
    signal MUX_787_wire : std_logic_vector(15 downto 0);
    signal MUX_794_wire : std_logic_vector(15 downto 0);
    signal MUX_817_wire : std_logic_vector(15 downto 0);
    signal MUX_870_wire : std_logic_vector(31 downto 0);
    signal MUX_871_wire : std_logic_vector(31 downto 0);
    signal MUX_880_wire : std_logic_vector(0 downto 0);
    signal MUX_886_wire : std_logic_vector(0 downto 0);
    signal MUX_893_wire : std_logic_vector(0 downto 0);
    signal MUX_899_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_801_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_822_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_830_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_838_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_846_wire : std_logic_vector(0 downto 0);
    signal OR_u16_u16_780_wire : std_logic_vector(15 downto 0);
    signal OR_u16_u16_795_wire : std_logic_vector(15 downto 0);
    signal OR_u1_u1_739_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_752_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_887_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_900_wire : std_logic_vector(0 downto 0);
    signal RPIPE_noblock_obuf_1_1_665_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_1_670_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_1_675_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_1_680_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_16_687_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_33_663_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_668_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_673_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_678_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_683_wire_constant : std_logic_vector(2 downto 0);
    signal SUB_u16_u16_811_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_815_wire : std_logic_vector(15 downto 0);
    signal active_packet_681 : std_logic_vector(2 downto 0);
    signal data_to_out_873 : std_logic_vector(31 downto 0);
    signal down_counter_685 : std_logic_vector(15 downto 0);
    signal konst_691_wire_constant : std_logic_vector(2 downto 0);
    signal konst_696_wire_constant : std_logic_vector(32 downto 0);
    signal konst_701_wire_constant : std_logic_vector(32 downto 0);
    signal konst_706_wire_constant : std_logic_vector(32 downto 0);
    signal konst_711_wire_constant : std_logic_vector(32 downto 0);
    signal konst_728_wire_constant : std_logic_vector(2 downto 0);
    signal konst_731_wire_constant : std_logic_vector(0 downto 0);
    signal konst_734_wire_constant : std_logic_vector(2 downto 0);
    signal konst_737_wire_constant : std_logic_vector(0 downto 0);
    signal konst_741_wire_constant : std_logic_vector(2 downto 0);
    signal konst_744_wire_constant : std_logic_vector(0 downto 0);
    signal konst_747_wire_constant : std_logic_vector(2 downto 0);
    signal konst_750_wire_constant : std_logic_vector(0 downto 0);
    signal konst_767_wire_constant : std_logic_vector(2 downto 0);
    signal konst_771_wire_constant : std_logic_vector(15 downto 0);
    signal konst_774_wire_constant : std_logic_vector(2 downto 0);
    signal konst_778_wire_constant : std_logic_vector(15 downto 0);
    signal konst_782_wire_constant : std_logic_vector(2 downto 0);
    signal konst_786_wire_constant : std_logic_vector(15 downto 0);
    signal konst_789_wire_constant : std_logic_vector(2 downto 0);
    signal konst_793_wire_constant : std_logic_vector(15 downto 0);
    signal konst_800_wire_constant : std_logic_vector(2 downto 0);
    signal konst_803_wire_constant : std_logic_vector(15 downto 0);
    signal konst_810_wire_constant : std_logic_vector(15 downto 0);
    signal konst_814_wire_constant : std_logic_vector(15 downto 0);
    signal konst_824_wire_constant : std_logic_vector(2 downto 0);
    signal konst_832_wire_constant : std_logic_vector(2 downto 0);
    signal konst_840_wire_constant : std_logic_vector(2 downto 0);
    signal konst_848_wire_constant : std_logic_vector(2 downto 0);
    signal konst_854_wire_constant : std_logic_vector(2 downto 0);
    signal konst_859_wire_constant : std_logic_vector(2 downto 0);
    signal konst_864_wire_constant : std_logic_vector(2 downto 0);
    signal konst_876_wire_constant : std_logic_vector(2 downto 0);
    signal konst_879_wire_constant : std_logic_vector(0 downto 0);
    signal konst_882_wire_constant : std_logic_vector(2 downto 0);
    signal konst_885_wire_constant : std_logic_vector(0 downto 0);
    signal konst_889_wire_constant : std_logic_vector(2 downto 0);
    signal konst_892_wire_constant : std_logic_vector(0 downto 0);
    signal konst_895_wire_constant : std_logic_vector(2 downto 0);
    signal konst_898_wire_constant : std_logic_vector(0 downto 0);
    signal konst_917_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_764 : std_logic_vector(2 downto 0);
    signal next_active_packet_764_684_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_819 : std_logic_vector(15 downto 0);
    signal next_down_counter_819_688_buffered : std_logic_vector(15 downto 0);
    signal next_pkt_with_priority_764 : std_logic_vector(2 downto 0);
    signal next_pkt_with_priority_764_692_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_698 : std_logic_vector(0 downto 0);
    signal p2_valid_703 : std_logic_vector(0 downto 0);
    signal p3_valid_708 : std_logic_vector(0 downto 0);
    signal p4_valid_713 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_661 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_666 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_671 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_676 : std_logic_vector(32 downto 0);
    signal pkt_with_priority_689 : std_logic_vector(2 downto 0);
    signal read_from_1_827 : std_logic_vector(0 downto 0);
    signal read_from_2_835 : std_logic_vector(0 downto 0);
    signal read_from_3_843 : std_logic_vector(0 downto 0);
    signal read_from_4_851 : std_logic_vector(0 downto 0);
    signal send_flag_902 : std_logic_vector(0 downto 0);
    signal slice_770_wire : std_logic_vector(15 downto 0);
    signal slice_777_wire : std_logic_vector(15 downto 0);
    signal slice_785_wire : std_logic_vector(15 downto 0);
    signal slice_792_wire : std_logic_vector(15 downto 0);
    signal slice_857_wire : std_logic_vector(31 downto 0);
    signal slice_862_wire : std_logic_vector(31 downto 0);
    signal slice_867_wire : std_logic_vector(31 downto 0);
    signal slice_869_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_806 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_length_797 : std_logic_vector(15 downto 0);
    signal valid_active_pkt_word_read_754 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_16_687_wire_constant <= "0000000000000000";
    R_ZERO_33_663_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_668_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_673_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_678_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_683_wire_constant <= "000";
    konst_691_wire_constant <= "001";
    konst_696_wire_constant <= "000000000000000000000000000100000";
    konst_701_wire_constant <= "000000000000000000000000000100000";
    konst_706_wire_constant <= "000000000000000000000000000100000";
    konst_711_wire_constant <= "000000000000000000000000000100000";
    konst_728_wire_constant <= "001";
    konst_731_wire_constant <= "0";
    konst_734_wire_constant <= "010";
    konst_737_wire_constant <= "0";
    konst_741_wire_constant <= "011";
    konst_744_wire_constant <= "0";
    konst_747_wire_constant <= "100";
    konst_750_wire_constant <= "0";
    konst_767_wire_constant <= "001";
    konst_771_wire_constant <= "0000000000000000";
    konst_774_wire_constant <= "010";
    konst_778_wire_constant <= "0000000000000000";
    konst_782_wire_constant <= "011";
    konst_786_wire_constant <= "0000000000000000";
    konst_789_wire_constant <= "100";
    konst_793_wire_constant <= "0000000000000000";
    konst_800_wire_constant <= "000";
    konst_803_wire_constant <= "0000000000000000";
    konst_810_wire_constant <= "0000000000000001";
    konst_814_wire_constant <= "0000000000000001";
    konst_824_wire_constant <= "001";
    konst_832_wire_constant <= "010";
    konst_840_wire_constant <= "011";
    konst_848_wire_constant <= "100";
    konst_854_wire_constant <= "001";
    konst_859_wire_constant <= "010";
    konst_864_wire_constant <= "011";
    konst_876_wire_constant <= "001";
    konst_879_wire_constant <= "0";
    konst_882_wire_constant <= "010";
    konst_885_wire_constant <= "0";
    konst_889_wire_constant <= "011";
    konst_892_wire_constant <= "0";
    konst_895_wire_constant <= "100";
    konst_898_wire_constant <= "0";
    konst_917_wire_constant <= "1";
    phi_stmt_661: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_663_wire_constant & RPIPE_noblock_obuf_1_1_665_wire;
      req <= phi_stmt_661_req_0 & phi_stmt_661_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_661",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_661_ack_0,
          idata => idata,
          odata => pkt_1_e_word_661,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_661
    phi_stmt_666: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_668_wire_constant & RPIPE_noblock_obuf_2_1_670_wire;
      req <= phi_stmt_666_req_0 & phi_stmt_666_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_666",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_666_ack_0,
          idata => idata,
          odata => pkt_2_e_word_666,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_666
    phi_stmt_671: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_673_wire_constant & RPIPE_noblock_obuf_3_1_675_wire;
      req <= phi_stmt_671_req_0 & phi_stmt_671_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_671",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_671_ack_0,
          idata => idata,
          odata => pkt_3_e_word_671,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_671
    phi_stmt_676: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_678_wire_constant & RPIPE_noblock_obuf_4_1_680_wire;
      req <= phi_stmt_676_req_0 & phi_stmt_676_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_676",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_676_ack_0,
          idata => idata,
          odata => pkt_4_e_word_676,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_676
    phi_stmt_681: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_683_wire_constant & next_active_packet_764_684_buffered;
      req <= phi_stmt_681_req_0 & phi_stmt_681_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_681",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_681_ack_0,
          idata => idata,
          odata => active_packet_681,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_681
    phi_stmt_685: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_16_687_wire_constant & next_down_counter_819_688_buffered;
      req <= phi_stmt_685_req_0 & phi_stmt_685_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_685",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_685_ack_0,
          idata => idata,
          odata => down_counter_685,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_685
    phi_stmt_689: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_691_wire_constant & next_pkt_with_priority_764_692_buffered;
      req <= phi_stmt_689_req_0 & phi_stmt_689_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_689",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_689_ack_0,
          idata => idata,
          odata => pkt_with_priority_689,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_689
    -- flow-through select operator MUX_732_inst
    MUX_732_wire <= p1_valid_698 when (EQ_u3_u1_729_wire(0) /=  '0') else konst_731_wire_constant;
    -- flow-through select operator MUX_738_inst
    MUX_738_wire <= p2_valid_703 when (EQ_u3_u1_735_wire(0) /=  '0') else konst_737_wire_constant;
    -- flow-through select operator MUX_745_inst
    MUX_745_wire <= p3_valid_708 when (EQ_u3_u1_742_wire(0) /=  '0') else konst_744_wire_constant;
    -- flow-through select operator MUX_751_inst
    MUX_751_wire <= p4_valid_713 when (EQ_u3_u1_748_wire(0) /=  '0') else konst_750_wire_constant;
    -- flow-through select operator MUX_772_inst
    MUX_772_wire <= slice_770_wire when (EQ_u3_u1_768_wire(0) /=  '0') else konst_771_wire_constant;
    -- flow-through select operator MUX_779_inst
    MUX_779_wire <= slice_777_wire when (EQ_u3_u1_775_wire(0) /=  '0') else konst_778_wire_constant;
    -- flow-through select operator MUX_787_inst
    MUX_787_wire <= slice_785_wire when (EQ_u3_u1_783_wire(0) /=  '0') else konst_786_wire_constant;
    -- flow-through select operator MUX_794_inst
    MUX_794_wire <= slice_792_wire when (EQ_u3_u1_790_wire(0) /=  '0') else konst_793_wire_constant;
    -- flow-through select operator MUX_817_inst
    MUX_817_wire <= SUB_u16_u16_815_wire when (valid_active_pkt_word_read_754(0) /=  '0') else down_counter_685;
    -- flow-through select operator MUX_818_inst
    next_down_counter_819 <= SUB_u16_u16_811_wire when (started_new_packet_806(0) /=  '0') else MUX_817_wire;
    -- flow-through select operator MUX_870_inst
    MUX_870_wire <= slice_867_wire when (EQ_u3_u1_865_wire(0) /=  '0') else slice_869_wire;
    -- flow-through select operator MUX_871_inst
    MUX_871_wire <= slice_862_wire when (EQ_u3_u1_860_wire(0) /=  '0') else MUX_870_wire;
    -- flow-through select operator MUX_872_inst
    data_to_out_873 <= slice_857_wire when (EQ_u3_u1_855_wire(0) /=  '0') else MUX_871_wire;
    -- flow-through select operator MUX_880_inst
    MUX_880_wire <= p1_valid_698 when (EQ_u3_u1_877_wire(0) /=  '0') else konst_879_wire_constant;
    -- flow-through select operator MUX_886_inst
    MUX_886_wire <= p2_valid_703 when (EQ_u3_u1_883_wire(0) /=  '0') else konst_885_wire_constant;
    -- flow-through select operator MUX_893_inst
    MUX_893_wire <= p3_valid_708 when (EQ_u3_u1_890_wire(0) /=  '0') else konst_892_wire_constant;
    -- flow-through select operator MUX_899_inst
    MUX_899_wire <= p4_valid_713 when (EQ_u3_u1_896_wire(0) /=  '0') else konst_898_wire_constant;
    -- flow-through slice operator slice_770_inst
    slice_770_wire <= pkt_1_e_word_661(23 downto 8);
    -- flow-through slice operator slice_777_inst
    slice_777_wire <= pkt_2_e_word_666(23 downto 8);
    -- flow-through slice operator slice_785_inst
    slice_785_wire <= pkt_3_e_word_671(23 downto 8);
    -- flow-through slice operator slice_792_inst
    slice_792_wire <= pkt_4_e_word_676(23 downto 8);
    -- flow-through slice operator slice_857_inst
    slice_857_wire <= pkt_1_e_word_661(31 downto 0);
    -- flow-through slice operator slice_862_inst
    slice_862_wire <= pkt_2_e_word_666(31 downto 0);
    -- flow-through slice operator slice_867_inst
    slice_867_wire <= pkt_3_e_word_671(31 downto 0);
    -- flow-through slice operator slice_869_inst
    slice_869_wire <= pkt_4_e_word_676(31 downto 0);
    next_active_packet_764_684_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_764_684_buf_req_0;
      next_active_packet_764_684_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_764_684_buf_req_1;
      next_active_packet_764_684_buf_ack_1<= rack(0);
      next_active_packet_764_684_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_764_684_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_764_684_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_819_688_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_819_688_buf_req_0;
      next_down_counter_819_688_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_819_688_buf_req_1;
      next_down_counter_819_688_buf_ack_1<= rack(0);
      next_down_counter_819_688_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_819_688_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_819_688_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_with_priority_764_692_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_with_priority_764_692_buf_req_0;
      next_pkt_with_priority_764_692_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_with_priority_764_692_buf_req_1;
      next_pkt_with_priority_764_692_buf_ack_1<= rack(0);
      next_pkt_with_priority_764_692_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_with_priority_764_692_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_with_priority_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_with_priority_764_692_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_659_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_917_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_659_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_659_branch_req_0,
          ack0 => do_while_stmt_659_branch_ack_0,
          ack1 => do_while_stmt_659_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_805_inst
    process(NEQ_u3_u1_801_wire, EQ_u16_u1_804_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u3_u1_801_wire, EQ_u16_u1_804_wire, tmp_var);
      started_new_packet_806 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_697_inst
    process(pkt_1_e_word_661) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_661, konst_696_wire_constant, tmp_var);
      p1_valid_698 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_702_inst
    process(pkt_2_e_word_666) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_666, konst_701_wire_constant, tmp_var);
      p2_valid_703 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_707_inst
    process(pkt_3_e_word_671) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_671, konst_706_wire_constant, tmp_var);
      p3_valid_708 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_712_inst
    process(pkt_4_e_word_676) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_676, konst_711_wire_constant, tmp_var);
      p4_valid_713 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_804_inst
    process(down_counter_685) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_685, konst_803_wire_constant, tmp_var);
      EQ_u16_u1_804_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_729_inst
    process(active_packet_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_681, konst_728_wire_constant, tmp_var);
      EQ_u3_u1_729_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_735_inst
    process(active_packet_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_681, konst_734_wire_constant, tmp_var);
      EQ_u3_u1_735_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_742_inst
    process(active_packet_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_681, konst_741_wire_constant, tmp_var);
      EQ_u3_u1_742_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_748_inst
    process(active_packet_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_681, konst_747_wire_constant, tmp_var);
      EQ_u3_u1_748_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_768_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_767_wire_constant, tmp_var);
      EQ_u3_u1_768_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_775_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_774_wire_constant, tmp_var);
      EQ_u3_u1_775_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_783_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_782_wire_constant, tmp_var);
      EQ_u3_u1_783_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_790_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_789_wire_constant, tmp_var);
      EQ_u3_u1_790_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_825_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_824_wire_constant, tmp_var);
      EQ_u3_u1_825_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_833_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_832_wire_constant, tmp_var);
      EQ_u3_u1_833_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_841_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_840_wire_constant, tmp_var);
      EQ_u3_u1_841_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_849_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_848_wire_constant, tmp_var);
      EQ_u3_u1_849_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_855_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_854_wire_constant, tmp_var);
      EQ_u3_u1_855_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_860_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_859_wire_constant, tmp_var);
      EQ_u3_u1_860_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_865_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_864_wire_constant, tmp_var);
      EQ_u3_u1_865_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_877_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_876_wire_constant, tmp_var);
      EQ_u3_u1_877_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_883_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_882_wire_constant, tmp_var);
      EQ_u3_u1_883_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_890_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_889_wire_constant, tmp_var);
      EQ_u3_u1_890_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_896_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_764, konst_895_wire_constant, tmp_var);
      EQ_u3_u1_896_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_801_inst
    process(next_active_packet_764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_764, konst_800_wire_constant, tmp_var);
      NEQ_u3_u1_801_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_822_inst
    process(p1_valid_698) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_698, tmp_var);
      NOT_u1_u1_822_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_830_inst
    process(p2_valid_703) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_703, tmp_var);
      NOT_u1_u1_830_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_838_inst
    process(p3_valid_708) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_708, tmp_var);
      NOT_u1_u1_838_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_846_inst
    process(p4_valid_713) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_713, tmp_var);
      NOT_u1_u1_846_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_780_inst
    process(MUX_772_wire, MUX_779_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_772_wire, MUX_779_wire, tmp_var);
      OR_u16_u16_780_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_795_inst
    process(MUX_787_wire, MUX_794_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_787_wire, MUX_794_wire, tmp_var);
      OR_u16_u16_795_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_796_inst
    process(OR_u16_u16_780_wire, OR_u16_u16_795_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u16_u16_780_wire, OR_u16_u16_795_wire, tmp_var);
      valid_active_pkt_length_797 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_739_inst
    process(MUX_732_wire, MUX_738_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_732_wire, MUX_738_wire, tmp_var);
      OR_u1_u1_739_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_752_inst
    process(MUX_745_wire, MUX_751_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_745_wire, MUX_751_wire, tmp_var);
      OR_u1_u1_752_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_753_inst
    process(OR_u1_u1_739_wire, OR_u1_u1_752_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_739_wire, OR_u1_u1_752_wire, tmp_var);
      valid_active_pkt_word_read_754 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_826_inst
    process(NOT_u1_u1_822_wire, EQ_u3_u1_825_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_822_wire, EQ_u3_u1_825_wire, tmp_var);
      read_from_1_827 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_834_inst
    process(NOT_u1_u1_830_wire, EQ_u3_u1_833_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_830_wire, EQ_u3_u1_833_wire, tmp_var);
      read_from_2_835 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_842_inst
    process(NOT_u1_u1_838_wire, EQ_u3_u1_841_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_838_wire, EQ_u3_u1_841_wire, tmp_var);
      read_from_3_843 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_850_inst
    process(NOT_u1_u1_846_wire, EQ_u3_u1_849_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_846_wire, EQ_u3_u1_849_wire, tmp_var);
      read_from_4_851 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_887_inst
    process(MUX_880_wire, MUX_886_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_880_wire, MUX_886_wire, tmp_var);
      OR_u1_u1_887_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_900_inst
    process(MUX_893_wire, MUX_899_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_893_wire, MUX_899_wire, tmp_var);
      OR_u1_u1_900_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_901_inst
    process(OR_u1_u1_887_wire, OR_u1_u1_900_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_887_wire, OR_u1_u1_900_wire, tmp_var);
      send_flag_902 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_811_inst
    process(valid_active_pkt_length_797) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(valid_active_pkt_length_797, konst_810_wire_constant, tmp_var);
      SUB_u16_u16_811_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_815_inst
    process(down_counter_685) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_685, konst_814_wire_constant, tmp_var);
      SUB_u16_u16_815_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_1_665_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_1_665_inst_req_0;
      RPIPE_noblock_obuf_1_1_665_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_1_665_inst_req_1;
      RPIPE_noblock_obuf_1_1_665_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_827(0);
      RPIPE_noblock_obuf_1_1_665_wire <= data_out(32 downto 0);
      noblock_obuf_1_1_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_1_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_1_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_1_pipe_read_req(0),
          oack => noblock_obuf_1_1_pipe_read_ack(0),
          odata => noblock_obuf_1_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_1_670_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_1_670_inst_req_0;
      RPIPE_noblock_obuf_2_1_670_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_1_670_inst_req_1;
      RPIPE_noblock_obuf_2_1_670_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_835(0);
      RPIPE_noblock_obuf_2_1_670_wire <= data_out(32 downto 0);
      noblock_obuf_2_1_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_1_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_1_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_1_pipe_read_req(0),
          oack => noblock_obuf_2_1_pipe_read_ack(0),
          odata => noblock_obuf_2_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_1_675_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_1_675_inst_req_0;
      RPIPE_noblock_obuf_3_1_675_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_1_675_inst_req_1;
      RPIPE_noblock_obuf_3_1_675_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_843(0);
      RPIPE_noblock_obuf_3_1_675_wire <= data_out(32 downto 0);
      noblock_obuf_3_1_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_1_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_1_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_1_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_1_pipe_read_req(0),
          oack => noblock_obuf_3_1_pipe_read_ack(0),
          odata => noblock_obuf_3_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_1_680_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_1_680_inst_req_0;
      RPIPE_noblock_obuf_4_1_680_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_1_680_inst_req_1;
      RPIPE_noblock_obuf_4_1_680_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_851(0);
      RPIPE_noblock_obuf_4_1_680_wire <= data_out(32 downto 0);
      noblock_obuf_4_1_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_1_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_1_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_1_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_1_pipe_read_req(0),
          oack => noblock_obuf_4_1_pipe_read_ack(0),
          odata => noblock_obuf_4_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_1_904_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_1_904_inst_req_0;
      WPIPE_out_data_1_904_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_1_904_inst_req_1;
      WPIPE_out_data_1_904_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_902(0);
      data_in <= data_to_out_873;
      out_data_1_write_0_gI: SplitGuardInterface generic map(name => "out_data_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_1_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_1", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_1_pipe_write_req(0),
          oack => out_data_1_pipe_write_ack(0),
          odata => out_data_1_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_1893: prioritySelect_Volatile port map(down_counter => down_counter_685, active_packet => active_packet_681, pkt_with_priority => pkt_with_priority_689, p1_valid => p1_valid_698, p2_valid => p2_valid_703, p3_valid => p3_valid_708, p4_valid => p4_valid_713, next_active_packet => next_active_packet_764, next_pkt_with_priority => next_pkt_with_priority_764); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_1_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_2_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_2_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_2_Daemon;
architecture outputPort_2_Daemon_arch of outputPort_2_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_2_Daemon_CP_1176_start: Boolean;
  signal outputPort_2_Daemon_CP_1176_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(15 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_with_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_with_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal next_down_counter_1082_951_buf_ack_1 : boolean;
  signal next_pkt_with_priority_1027_955_buf_ack_1 : boolean;
  signal WPIPE_out_data_2_1167_inst_ack_0 : boolean;
  signal next_pkt_with_priority_1027_955_buf_req_1 : boolean;
  signal WPIPE_out_data_2_1167_inst_req_0 : boolean;
  signal next_down_counter_1082_951_buf_ack_0 : boolean;
  signal next_down_counter_1082_951_buf_req_0 : boolean;
  signal WPIPE_out_data_2_1167_inst_req_1 : boolean;
  signal phi_stmt_952_req_0 : boolean;
  signal WPIPE_out_data_2_1167_inst_ack_1 : boolean;
  signal next_down_counter_1082_951_buf_req_1 : boolean;
  signal phi_stmt_948_ack_0 : boolean;
  signal next_pkt_with_priority_1027_955_buf_req_0 : boolean;
  signal phi_stmt_952_req_1 : boolean;
  signal next_pkt_with_priority_1027_955_buf_ack_0 : boolean;
  signal do_while_stmt_922_branch_req_0 : boolean;
  signal phi_stmt_924_req_1 : boolean;
  signal phi_stmt_948_req_1 : boolean;
  signal phi_stmt_952_ack_0 : boolean;
  signal phi_stmt_948_req_0 : boolean;
  signal do_while_stmt_922_branch_ack_0 : boolean;
  signal phi_stmt_924_req_0 : boolean;
  signal phi_stmt_924_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_928_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_928_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_928_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_2_928_inst_ack_1 : boolean;
  signal phi_stmt_929_req_1 : boolean;
  signal phi_stmt_929_req_0 : boolean;
  signal phi_stmt_929_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_933_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_933_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_933_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_2_933_inst_ack_1 : boolean;
  signal do_while_stmt_922_branch_ack_1 : boolean;
  signal phi_stmt_934_req_1 : boolean;
  signal phi_stmt_934_req_0 : boolean;
  signal phi_stmt_934_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_938_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_938_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_938_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_2_938_inst_ack_1 : boolean;
  signal phi_stmt_939_req_1 : boolean;
  signal phi_stmt_939_req_0 : boolean;
  signal phi_stmt_939_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_943_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_943_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_943_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_2_943_inst_ack_1 : boolean;
  signal phi_stmt_944_req_1 : boolean;
  signal phi_stmt_944_req_0 : boolean;
  signal phi_stmt_944_ack_0 : boolean;
  signal next_active_packet_1027_947_buf_req_0 : boolean;
  signal next_active_packet_1027_947_buf_ack_0 : boolean;
  signal next_active_packet_1027_947_buf_req_1 : boolean;
  signal next_active_packet_1027_947_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_2_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_2_Daemon_CP_1176_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_2_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_2_Daemon_CP_1176: Block -- control-path 
    signal outputPort_2_Daemon_CP_1176_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_2_Daemon_CP_1176_elements(0) <= outputPort_2_Daemon_CP_1176_start;
    outputPort_2_Daemon_CP_1176_symbol <= outputPort_2_Daemon_CP_1176_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_921/$entry
      -- CP-element group 0: 	 branch_block_stmt_921/do_while_stmt_922__entry__
      -- CP-element group 0: 	 branch_block_stmt_921/branch_block_stmt_921__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_921/do_while_stmt_922__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_921/$exit
      -- CP-element group 1: 	 branch_block_stmt_921/branch_block_stmt_921__exit__
      -- 
    outputPort_2_Daemon_CP_1176_elements(1) <= outputPort_2_Daemon_CP_1176_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_921/do_while_stmt_922/$entry
      -- CP-element group 2: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922__entry__
      -- 
    outputPort_2_Daemon_CP_1176_elements(2) <= outputPort_2_Daemon_CP_1176_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922__exit__
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_921/do_while_stmt_922/loop_back
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	159 
    -- CP-element group 5: 	160 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_921/do_while_stmt_922/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_921/do_while_stmt_922/condition_done
      -- CP-element group 5: 	 branch_block_stmt_921/do_while_stmt_922/loop_taken/$entry
      -- 
    outputPort_2_Daemon_CP_1176_elements(5) <= outputPort_2_Daemon_CP_1176_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_921/do_while_stmt_922/loop_body_done
      -- 
    outputPort_2_Daemon_CP_1176_elements(6) <= outputPort_2_Daemon_CP_1176_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	104 
    -- CP-element group 7: 	83 
    -- CP-element group 7: 	122 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	42 
    -- CP-element group 7: 	63 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/back_edge_to_loop_body
      -- 
    outputPort_2_Daemon_CP_1176_elements(7) <= outputPort_2_Daemon_CP_1176_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	85 
    -- CP-element group 8: 	124 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	44 
    -- CP-element group 8: 	106 
    -- CP-element group 8: 	65 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/first_time_through_loop_body
      -- 
    outputPort_2_Daemon_CP_1176_elements(8) <= outputPort_2_Daemon_CP_1176_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	99 
    -- CP-element group 9: 	79 
    -- CP-element group 9: 	117 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	135 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	57 
    -- CP-element group 9: 	58 
    -- CP-element group 9: 	78 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/loop_body_start
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/condition_evaluated
      -- 
    condition_evaluated_1200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(10), ack => do_while_stmt_922_branch_req_0); -- 
    outputPort_2_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(157) & outputPort_2_Daemon_CP_1176_elements(14);
      gj_outputPort_2_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	117 
    -- CP-element group 11: 	135 
    -- CP-element group 11: 	98 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	100 
    -- CP-element group 11: 	119 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	38 
    -- CP-element group 11: 	59 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_sample_start__ps
      -- 
    outputPort_2_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(117) & outputPort_2_Daemon_CP_1176_elements(135) & outputPort_2_Daemon_CP_1176_elements(98) & outputPort_2_Daemon_CP_1176_elements(15) & outputPort_2_Daemon_CP_1176_elements(36) & outputPort_2_Daemon_CP_1176_elements(57) & outputPort_2_Daemon_CP_1176_elements(78) & outputPort_2_Daemon_CP_1176_elements(14);
      gj_outputPort_2_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	120 
    -- CP-element group 12: 	80 
    -- CP-element group 12: 	101 
    -- CP-element group 12: 	138 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	39 
    -- CP-element group 12: 	60 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	117 
    -- CP-element group 12: 	135 
    -- CP-element group 12: 	98 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	57 
    -- CP-element group 12: 	78 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_sample_completed_
      -- 
    outputPort_2_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(120) & outputPort_2_Daemon_CP_1176_elements(80) & outputPort_2_Daemon_CP_1176_elements(101) & outputPort_2_Daemon_CP_1176_elements(138) & outputPort_2_Daemon_CP_1176_elements(18) & outputPort_2_Daemon_CP_1176_elements(39) & outputPort_2_Daemon_CP_1176_elements(60);
      gj_outputPort_2_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	136 
    -- CP-element group 13: 	99 
    -- CP-element group 13: 	79 
    -- CP-element group 13: 	118 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	58 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	81 
    -- CP-element group 13: 	102 
    -- CP-element group 13: 	139 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	40 
    -- CP-element group 13: 	61 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/aggregated_phi_update_req
      -- 
    outputPort_2_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(136) & outputPort_2_Daemon_CP_1176_elements(99) & outputPort_2_Daemon_CP_1176_elements(79) & outputPort_2_Daemon_CP_1176_elements(118) & outputPort_2_Daemon_CP_1176_elements(16) & outputPort_2_Daemon_CP_1176_elements(37) & outputPort_2_Daemon_CP_1176_elements(58);
      gj_outputPort_2_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	121 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	82 
    -- CP-element group 14: 	103 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	41 
    -- CP-element group 14: 	62 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_2_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(121) & outputPort_2_Daemon_CP_1176_elements(140) & outputPort_2_Daemon_CP_1176_elements(82) & outputPort_2_Daemon_CP_1176_elements(103) & outputPort_2_Daemon_CP_1176_elements(20) & outputPort_2_Daemon_CP_1176_elements(41) & outputPort_2_Daemon_CP_1176_elements(62);
      gj_outputPort_2_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(17) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(19) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(21) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_loopback_sample_req_ps
      -- 
    phi_stmt_924_loopback_sample_req_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_924_loopback_sample_req_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(22), ack => phi_stmt_924_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(23) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_entry_sample_req_ps
      -- 
    phi_stmt_924_entry_sample_req_1218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_924_entry_sample_req_1218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(24), ack => phi_stmt_924_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_924_phi_mux_ack_ps
      -- 
    phi_stmt_924_phi_mux_ack_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_924_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_926_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_926_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_926_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_926_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_926_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_926_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_926_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(28) <= outputPort_2_Daemon_CP_1176_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_926_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(27), ack => outputPort_2_Daemon_CP_1176_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	35 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_Sample/rr
      -- 
    rr_1242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(32), ack => RPIPE_noblock_obuf_1_2_928_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(30) & outputPort_2_Daemon_CP_1176_elements(35);
      gj_outputPort_2_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: 	34 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_update_start_
      -- CP-element group 33: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_Update/cr
      -- 
    cr_1247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(33), ack => RPIPE_noblock_obuf_1_2_928_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(31) & outputPort_2_Daemon_CP_1176_elements(34);
      gj_outputPort_2_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	33 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_Sample/ra
      -- 
    ra_1243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_2_928_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	32 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_1_2_928_Update/ca
      -- 
    ca_1248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_2_928_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	11 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	155 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	11 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(38) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	12 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	13 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(40) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	154 
    -- CP-element group 41: 	14 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	7 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(42) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_loopback_sample_req_ps
      -- 
    phi_stmt_929_loopback_sample_req_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_929_loopback_sample_req_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(43), ack => phi_stmt_929_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	8 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(44) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_entry_sample_req
      -- CP-element group 45: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_entry_sample_req_ps
      -- 
    phi_stmt_929_entry_sample_req_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_929_entry_sample_req_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(45), ack => phi_stmt_929_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_929_phi_mux_ack_ps
      -- 
    phi_stmt_929_phi_mux_ack_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_929_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_931_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_931_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_931_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_931_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_931_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_931_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_931_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(49) <= outputPort_2_Daemon_CP_1176_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_931_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(48), ack => outputPort_2_Daemon_CP_1176_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_Sample/rr
      -- 
    rr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(53), ack => RPIPE_noblock_obuf_2_2_933_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(51) & outputPort_2_Daemon_CP_1176_elements(56);
      gj_outputPort_2_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: 	55 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_update_start_
      -- CP-element group 54: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_Update/cr
      -- 
    cr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(54), ack => RPIPE_noblock_obuf_2_2_933_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(52) & outputPort_2_Daemon_CP_1176_elements(55);
      gj_outputPort_2_Daemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	54 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_Sample/ra
      -- 
    ra_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_2_933_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_2_2_933_Update/ca
      -- 
    ca_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_2_933_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(56)); -- 
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	9 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	12 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	11 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	9 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	155 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	13 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	11 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(59) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	12 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	13 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(61) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	154 
    -- CP-element group 62: 	14 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	7 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(63) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_loopback_sample_req
      -- CP-element group 64: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_loopback_sample_req_ps
      -- 
    phi_stmt_934_loopback_sample_req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_934_loopback_sample_req_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(64), ack => phi_stmt_934_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	8 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(65) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_entry_sample_req
      -- CP-element group 66: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_entry_sample_req_ps
      -- 
    phi_stmt_934_entry_sample_req_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_934_entry_sample_req_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(66), ack => phi_stmt_934_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_phi_mux_ack
      -- CP-element group 67: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_934_phi_mux_ack_ps
      -- 
    phi_stmt_934_phi_mux_ack_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_934_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_936_sample_start__ps
      -- CP-element group 68: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_936_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_936_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_936_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_936_update_start__ps
      -- CP-element group 69: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_936_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_936_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(70) <= outputPort_2_Daemon_CP_1176_elements(71);
    -- CP-element group 71:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	70 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_936_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(69), ack => outputPort_2_Daemon_CP_1176_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	77 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_Sample/rr
      -- 
    rr_1330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(74), ack => RPIPE_noblock_obuf_3_2_938_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(72) & outputPort_2_Daemon_CP_1176_elements(77);
      gj_outputPort_2_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	76 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_update_start_
      -- CP-element group 75: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_Update/cr
      -- 
    cr_1335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(75), ack => RPIPE_noblock_obuf_3_2_938_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(73) & outputPort_2_Daemon_CP_1176_elements(76);
      gj_outputPort_2_Daemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	75 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_Sample/ra
      -- 
    ra_1331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_2_938_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(76)); -- 
    -- CP-element group 77:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	74 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_3_2_938_Update/ca
      -- 
    ca_1336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_2_938_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	12 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	11 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	9 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	155 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	13 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	12 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(80) is bound as output of CP function.
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	13 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(81) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	154 
    -- CP-element group 82: 	14 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(82) is bound as output of CP function.
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	7 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(83) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 84:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_loopback_sample_req
      -- CP-element group 84: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_loopback_sample_req_ps
      -- 
    phi_stmt_939_loopback_sample_req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_939_loopback_sample_req_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(84), ack => phi_stmt_939_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(84) is bound as output of CP function.
    -- CP-element group 85:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(85) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 86:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_entry_sample_req
      -- CP-element group 86: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_entry_sample_req_ps
      -- 
    phi_stmt_939_entry_sample_req_1350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_939_entry_sample_req_1350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(86), ack => phi_stmt_939_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_phi_mux_ack
      -- CP-element group 87: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_939_phi_mux_ack_ps
      -- 
    phi_stmt_939_phi_mux_ack_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_939_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_941_sample_start__ps
      -- CP-element group 88: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_941_sample_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_941_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_941_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_941_update_start__ps
      -- CP-element group 89: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_941_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_941_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(90) <= outputPort_2_Daemon_CP_1176_elements(91);
    -- CP-element group 91:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	90 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_33_941_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(89), ack => outputPort_2_Daemon_CP_1176_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	97 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_Sample/rr
      -- 
    rr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(94), ack => RPIPE_noblock_obuf_4_2_943_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(92) & outputPort_2_Daemon_CP_1176_elements(97);
      gj_outputPort_2_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_update_start_
      -- CP-element group 95: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_Update/cr
      -- 
    cr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(95), ack => RPIPE_noblock_obuf_4_2_943_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(96) & outputPort_2_Daemon_CP_1176_elements(93);
      gj_outputPort_2_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	95 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_sample_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_Sample/ra
      -- 
    ra_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_2_943_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	94 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_update_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/RPIPE_noblock_obuf_4_2_943_Update/ca
      -- 
    ca_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_2_943_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(97)); -- 
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	12 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	11 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	9 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	155 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	13 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	11 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(100) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 101:  join  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	12 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	13 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(102) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	154 
    -- CP-element group 103: 	14 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(103) is bound as output of CP function.
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	7 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(104) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 105:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_loopback_sample_req
      -- CP-element group 105: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_loopback_sample_req_ps
      -- 
    phi_stmt_944_loopback_sample_req_1391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_944_loopback_sample_req_1391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(105), ack => phi_stmt_944_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	8 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(106) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 107:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_entry_sample_req
      -- CP-element group 107: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_entry_sample_req_ps
      -- 
    phi_stmt_944_entry_sample_req_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_944_entry_sample_req_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(107), ack => phi_stmt_944_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_phi_mux_ack
      -- CP-element group 108: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_944_phi_mux_ack_ps
      -- 
    phi_stmt_944_phi_mux_ack_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_944_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(108)); -- 
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_3_946_sample_start__ps
      -- CP-element group 109: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_3_946_sample_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_3_946_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_3_946_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_3_946_update_start__ps
      -- CP-element group 110: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_3_946_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_3_946_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(111) <= outputPort_2_Daemon_CP_1176_elements(112);
    -- CP-element group 112:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	111 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_3_946_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(110), ack => outputPort_2_Daemon_CP_1176_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_sample_start__ps
      -- CP-element group 113: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_Sample/req
      -- 
    req_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(113), ack => next_active_packet_1027_947_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_update_start__ps
      -- CP-element group 114: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_update_start_
      -- CP-element group 114: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_Update/req
      -- 
    req_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(114), ack => next_active_packet_1027_947_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_sample_completed__ps
      -- CP-element group 115: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_Sample/ack
      -- 
    ack_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1027_947_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(115)); -- 
    -- CP-element group 116:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_update_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_active_packet_947_Update/ack
      -- 
    ack_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1027_947_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(116)); -- 
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	9 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	12 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	11 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	155 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	13 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	11 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(119) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	12 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(120) is bound as output of CP function.
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	154 
    -- CP-element group 121: 	14 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	7 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(122) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_loopback_sample_req_ps
      -- CP-element group 123: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_loopback_sample_req
      -- 
    phi_stmt_948_loopback_sample_req_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_948_loopback_sample_req_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(123), ack => phi_stmt_948_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(124) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_entry_sample_req_ps
      -- CP-element group 125: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_entry_sample_req
      -- 
    phi_stmt_948_entry_sample_req_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_948_entry_sample_req_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(125), ack => phi_stmt_948_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_phi_mux_ack
      -- CP-element group 126: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_948_phi_mux_ack_ps
      -- 
    phi_stmt_948_phi_mux_ack_1441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_948_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_16_950_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_16_950_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_16_950_sample_start__ps
      -- CP-element group 127: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_16_950_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_16_950_update_start_
      -- CP-element group 128: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_16_950_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_16_950_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(129) <= outputPort_2_Daemon_CP_1176_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_ZERO_16_950_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(128), ack => outputPort_2_Daemon_CP_1176_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_Sample/req
      -- CP-element group 131: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_sample_start__ps
      -- 
    req_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(131), ack => next_down_counter_1082_951_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_update_start_
      -- CP-element group 132: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_Update/req
      -- CP-element group 132: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_update_start__ps
      -- CP-element group 132: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_Update/$entry
      -- 
    req_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(132), ack => next_down_counter_1082_951_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_Sample/ack
      -- CP-element group 133: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_Sample/$exit
      -- 
    ack_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1082_951_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(133)); -- 
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_Update/ack
      -- CP-element group 134: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_down_counter_951_update_completed_
      -- 
    ack_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1082_951_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	9 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	11 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	155 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	13 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(137) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	12 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	13 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(139) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_update_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(141) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_loopback_sample_req_ps
      -- 
    phi_stmt_952_loopback_sample_req_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_952_loopback_sample_req_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(142), ack => phi_stmt_952_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(143) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_entry_sample_req_ps
      -- 
    phi_stmt_952_entry_sample_req_1482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_952_entry_sample_req_1482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(144), ack => phi_stmt_952_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_phi_mux_ack_ps
      -- CP-element group 145: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/phi_stmt_952_phi_mux_ack
      -- 
    phi_stmt_952_phi_mux_ack_1485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_952_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/konst_954_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/konst_954_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/konst_954_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/konst_954_sample_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/konst_954_update_start_
      -- CP-element group 147: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/konst_954_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/konst_954_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(148) <= outputPort_2_Daemon_CP_1176_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/konst_954_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(147), ack => outputPort_2_Daemon_CP_1176_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_sample_start__ps
      -- 
    req_1506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(150), ack => next_pkt_with_priority_1027_955_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_Update/req
      -- CP-element group 151: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_update_start_
      -- CP-element group 151: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_Update/$entry
      -- 
    req_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(151), ack => next_pkt_with_priority_1027_955_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_sample_completed_
      -- 
    ack_1507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_with_priority_1027_955_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/R_next_pkt_with_priority_955_update_completed_
      -- 
    ack_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_with_priority_1027_955_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	121 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	82 
    -- CP-element group 154: 	103 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	41 
    -- CP-element group 154: 	62 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_Sample/req
      -- CP-element group 154: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_sample_start_
      -- 
    req_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(154), ack => WPIPE_out_data_2_1167_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(121) & outputPort_2_Daemon_CP_1176_elements(140) & outputPort_2_Daemon_CP_1176_elements(82) & outputPort_2_Daemon_CP_1176_elements(103) & outputPort_2_Daemon_CP_1176_elements(20) & outputPort_2_Daemon_CP_1176_elements(41) & outputPort_2_Daemon_CP_1176_elements(62) & outputPort_2_Daemon_CP_1176_elements(156);
      gj_outputPort_2_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	136 
    -- CP-element group 155: 	99 
    -- CP-element group 155: 	79 
    -- CP-element group 155: 	118 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	37 
    -- CP-element group 155: 	58 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_Update/req
      -- CP-element group 155: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_update_start_
      -- CP-element group 155: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_sample_completed_
      -- 
    ack_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_2_1167_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(155)); -- 
    req_1526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(155), ack => WPIPE_out_data_2_1167_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/WPIPE_out_data_2_1167_Update/ack
      -- 
    ack_1527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_2_1167_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(9), ack => outputPort_2_Daemon_CP_1176_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_921/do_while_stmt_922/do_while_stmt_922_loop_body/$exit
      -- 
    outputPort_2_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(156) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_921/do_while_stmt_922/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_921/do_while_stmt_922/loop_exit/ack
      -- 
    ack_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_922_branch_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_921/do_while_stmt_922/loop_taken/$exit
      -- CP-element group 160: 	 branch_block_stmt_921/do_while_stmt_922/loop_taken/ack
      -- 
    ack_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_922_branch_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_921/do_while_stmt_922/$exit
      -- 
    outputPort_2_Daemon_CP_1176_elements(161) <= outputPort_2_Daemon_CP_1176_elements(3);
    outputPort_2_Daemon_do_while_stmt_922_terminator_1537: loop_terminator -- 
      generic map (name => " outputPort_2_Daemon_do_while_stmt_922_terminator_1537", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_2_Daemon_CP_1176_elements(6),loop_continue => outputPort_2_Daemon_CP_1176_elements(160),loop_terminate => outputPort_2_Daemon_CP_1176_elements(159),loop_back => outputPort_2_Daemon_CP_1176_elements(4),loop_exit => outputPort_2_Daemon_CP_1176_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_924_phi_seq_1249_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(23);
      outputPort_2_Daemon_CP_1176_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(26);
      outputPort_2_Daemon_CP_1176_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(28);
      outputPort_2_Daemon_CP_1176_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(21);
      outputPort_2_Daemon_CP_1176_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(34);
      outputPort_2_Daemon_CP_1176_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(35);
      outputPort_2_Daemon_CP_1176_elements(22) <= phi_mux_reqs(1);
      phi_stmt_924_phi_seq_1249 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_924_phi_seq_1249") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(17), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(18), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(19), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(20), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_929_phi_seq_1293_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(44);
      outputPort_2_Daemon_CP_1176_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(47);
      outputPort_2_Daemon_CP_1176_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(49);
      outputPort_2_Daemon_CP_1176_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(42);
      outputPort_2_Daemon_CP_1176_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(55);
      outputPort_2_Daemon_CP_1176_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(56);
      outputPort_2_Daemon_CP_1176_elements(43) <= phi_mux_reqs(1);
      phi_stmt_929_phi_seq_1293 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_929_phi_seq_1293") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(38), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(39), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(40), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(41), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_934_phi_seq_1337_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(65);
      outputPort_2_Daemon_CP_1176_elements(68)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(68);
      outputPort_2_Daemon_CP_1176_elements(69)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(70);
      outputPort_2_Daemon_CP_1176_elements(66) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(63);
      outputPort_2_Daemon_CP_1176_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(76);
      outputPort_2_Daemon_CP_1176_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(77);
      outputPort_2_Daemon_CP_1176_elements(64) <= phi_mux_reqs(1);
      phi_stmt_934_phi_seq_1337 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_934_phi_seq_1337") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(59), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(60), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(61), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(62), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(67), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_939_phi_seq_1381_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(85);
      outputPort_2_Daemon_CP_1176_elements(88)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(88);
      outputPort_2_Daemon_CP_1176_elements(89)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(90);
      outputPort_2_Daemon_CP_1176_elements(86) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(83);
      outputPort_2_Daemon_CP_1176_elements(92)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(96);
      outputPort_2_Daemon_CP_1176_elements(93)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(97);
      outputPort_2_Daemon_CP_1176_elements(84) <= phi_mux_reqs(1);
      phi_stmt_939_phi_seq_1381 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_939_phi_seq_1381") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(11), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(80), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(81), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(82), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(87), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_944_phi_seq_1425_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(106);
      outputPort_2_Daemon_CP_1176_elements(109)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(109);
      outputPort_2_Daemon_CP_1176_elements(110)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(111);
      outputPort_2_Daemon_CP_1176_elements(107) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(104);
      outputPort_2_Daemon_CP_1176_elements(113)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(115);
      outputPort_2_Daemon_CP_1176_elements(114)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(116);
      outputPort_2_Daemon_CP_1176_elements(105) <= phi_mux_reqs(1);
      phi_stmt_944_phi_seq_1425 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_944_phi_seq_1425") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(100), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(101), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(102), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(103), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(108), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_948_phi_seq_1469_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(124);
      outputPort_2_Daemon_CP_1176_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(127);
      outputPort_2_Daemon_CP_1176_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(129);
      outputPort_2_Daemon_CP_1176_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(122);
      outputPort_2_Daemon_CP_1176_elements(131)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(133);
      outputPort_2_Daemon_CP_1176_elements(132)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(134);
      outputPort_2_Daemon_CP_1176_elements(123) <= phi_mux_reqs(1);
      phi_stmt_948_phi_seq_1469 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_948_phi_seq_1469") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(119), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(120), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(13), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(121), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_952_phi_seq_1513_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(143);
      outputPort_2_Daemon_CP_1176_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(146);
      outputPort_2_Daemon_CP_1176_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(148);
      outputPort_2_Daemon_CP_1176_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(141);
      outputPort_2_Daemon_CP_1176_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(152);
      outputPort_2_Daemon_CP_1176_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(153);
      outputPort_2_Daemon_CP_1176_elements(142) <= phi_mux_reqs(1);
      phi_stmt_952_phi_seq_1513 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_952_phi_seq_1513") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(137), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(138), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(139), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(140), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1201_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_2_Daemon_CP_1176_elements(7);
        preds(1)  <= outputPort_2_Daemon_CP_1176_elements(8);
        entry_tmerge_1201 : transition_merge -- 
          generic map(name => " entry_tmerge_1201")
          port map (preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u16_u1_1067_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1005_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1011_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1031_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1038_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1046_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1053_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1088_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1096_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1104_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1112_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1118_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1123_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1128_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1140_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1146_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1153_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1159_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_992_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_998_wire : std_logic_vector(0 downto 0);
    signal MUX_1001_wire : std_logic_vector(0 downto 0);
    signal MUX_1008_wire : std_logic_vector(0 downto 0);
    signal MUX_1014_wire : std_logic_vector(0 downto 0);
    signal MUX_1035_wire : std_logic_vector(15 downto 0);
    signal MUX_1042_wire : std_logic_vector(15 downto 0);
    signal MUX_1050_wire : std_logic_vector(15 downto 0);
    signal MUX_1057_wire : std_logic_vector(15 downto 0);
    signal MUX_1080_wire : std_logic_vector(15 downto 0);
    signal MUX_1133_wire : std_logic_vector(31 downto 0);
    signal MUX_1134_wire : std_logic_vector(31 downto 0);
    signal MUX_1143_wire : std_logic_vector(0 downto 0);
    signal MUX_1149_wire : std_logic_vector(0 downto 0);
    signal MUX_1156_wire : std_logic_vector(0 downto 0);
    signal MUX_1162_wire : std_logic_vector(0 downto 0);
    signal MUX_995_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_1064_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1085_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1093_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1101_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1109_wire : std_logic_vector(0 downto 0);
    signal OR_u16_u16_1043_wire : std_logic_vector(15 downto 0);
    signal OR_u16_u16_1058_wire : std_logic_vector(15 downto 0);
    signal OR_u1_u1_1002_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1015_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1150_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1163_wire : std_logic_vector(0 downto 0);
    signal RPIPE_noblock_obuf_1_2_928_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_2_933_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_2_938_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_2_943_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_16_950_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_33_926_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_931_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_936_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_941_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_946_wire_constant : std_logic_vector(2 downto 0);
    signal SUB_u16_u16_1074_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_1078_wire : std_logic_vector(15 downto 0);
    signal active_packet_944 : std_logic_vector(2 downto 0);
    signal data_to_out_1136 : std_logic_vector(31 downto 0);
    signal down_counter_948 : std_logic_vector(15 downto 0);
    signal konst_1000_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1004_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1007_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1010_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1013_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1030_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1034_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1037_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1041_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1045_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1049_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1052_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1056_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1063_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1066_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1073_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1077_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1087_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1095_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1103_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1111_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1117_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1122_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1127_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1139_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1142_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1145_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1148_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1152_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1155_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1158_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1161_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1180_wire_constant : std_logic_vector(0 downto 0);
    signal konst_954_wire_constant : std_logic_vector(2 downto 0);
    signal konst_959_wire_constant : std_logic_vector(32 downto 0);
    signal konst_964_wire_constant : std_logic_vector(32 downto 0);
    signal konst_969_wire_constant : std_logic_vector(32 downto 0);
    signal konst_974_wire_constant : std_logic_vector(32 downto 0);
    signal konst_991_wire_constant : std_logic_vector(2 downto 0);
    signal konst_994_wire_constant : std_logic_vector(0 downto 0);
    signal konst_997_wire_constant : std_logic_vector(2 downto 0);
    signal next_active_packet_1027 : std_logic_vector(2 downto 0);
    signal next_active_packet_1027_947_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_1082 : std_logic_vector(15 downto 0);
    signal next_down_counter_1082_951_buffered : std_logic_vector(15 downto 0);
    signal next_pkt_with_priority_1027 : std_logic_vector(2 downto 0);
    signal next_pkt_with_priority_1027_955_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_961 : std_logic_vector(0 downto 0);
    signal p2_valid_966 : std_logic_vector(0 downto 0);
    signal p3_valid_971 : std_logic_vector(0 downto 0);
    signal p4_valid_976 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_924 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_929 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_934 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_939 : std_logic_vector(32 downto 0);
    signal pkt_with_priority_952 : std_logic_vector(2 downto 0);
    signal read_from_1_1090 : std_logic_vector(0 downto 0);
    signal read_from_2_1098 : std_logic_vector(0 downto 0);
    signal read_from_3_1106 : std_logic_vector(0 downto 0);
    signal read_from_4_1114 : std_logic_vector(0 downto 0);
    signal send_flag_1165 : std_logic_vector(0 downto 0);
    signal slice_1033_wire : std_logic_vector(15 downto 0);
    signal slice_1040_wire : std_logic_vector(15 downto 0);
    signal slice_1048_wire : std_logic_vector(15 downto 0);
    signal slice_1055_wire : std_logic_vector(15 downto 0);
    signal slice_1120_wire : std_logic_vector(31 downto 0);
    signal slice_1125_wire : std_logic_vector(31 downto 0);
    signal slice_1130_wire : std_logic_vector(31 downto 0);
    signal slice_1132_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1069 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_length_1060 : std_logic_vector(15 downto 0);
    signal valid_active_pkt_word_read_1017 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_16_950_wire_constant <= "0000000000000000";
    R_ZERO_33_926_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_931_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_936_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_941_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_946_wire_constant <= "000";
    konst_1000_wire_constant <= "0";
    konst_1004_wire_constant <= "011";
    konst_1007_wire_constant <= "0";
    konst_1010_wire_constant <= "100";
    konst_1013_wire_constant <= "0";
    konst_1030_wire_constant <= "001";
    konst_1034_wire_constant <= "0000000000000000";
    konst_1037_wire_constant <= "010";
    konst_1041_wire_constant <= "0000000000000000";
    konst_1045_wire_constant <= "011";
    konst_1049_wire_constant <= "0000000000000000";
    konst_1052_wire_constant <= "100";
    konst_1056_wire_constant <= "0000000000000000";
    konst_1063_wire_constant <= "000";
    konst_1066_wire_constant <= "0000000000000000";
    konst_1073_wire_constant <= "0000000000000001";
    konst_1077_wire_constant <= "0000000000000001";
    konst_1087_wire_constant <= "001";
    konst_1095_wire_constant <= "010";
    konst_1103_wire_constant <= "011";
    konst_1111_wire_constant <= "100";
    konst_1117_wire_constant <= "001";
    konst_1122_wire_constant <= "010";
    konst_1127_wire_constant <= "011";
    konst_1139_wire_constant <= "001";
    konst_1142_wire_constant <= "0";
    konst_1145_wire_constant <= "010";
    konst_1148_wire_constant <= "0";
    konst_1152_wire_constant <= "011";
    konst_1155_wire_constant <= "0";
    konst_1158_wire_constant <= "100";
    konst_1161_wire_constant <= "0";
    konst_1180_wire_constant <= "1";
    konst_954_wire_constant <= "001";
    konst_959_wire_constant <= "000000000000000000000000000100000";
    konst_964_wire_constant <= "000000000000000000000000000100000";
    konst_969_wire_constant <= "000000000000000000000000000100000";
    konst_974_wire_constant <= "000000000000000000000000000100000";
    konst_991_wire_constant <= "001";
    konst_994_wire_constant <= "0";
    konst_997_wire_constant <= "010";
    phi_stmt_924: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_926_wire_constant & RPIPE_noblock_obuf_1_2_928_wire;
      req <= phi_stmt_924_req_0 & phi_stmt_924_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_924",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_924_ack_0,
          idata => idata,
          odata => pkt_1_e_word_924,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_924
    phi_stmt_929: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_931_wire_constant & RPIPE_noblock_obuf_2_2_933_wire;
      req <= phi_stmt_929_req_0 & phi_stmt_929_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_929",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_929_ack_0,
          idata => idata,
          odata => pkt_2_e_word_929,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_929
    phi_stmt_934: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_936_wire_constant & RPIPE_noblock_obuf_3_2_938_wire;
      req <= phi_stmt_934_req_0 & phi_stmt_934_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_934",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_934_ack_0,
          idata => idata,
          odata => pkt_3_e_word_934,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_934
    phi_stmt_939: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_941_wire_constant & RPIPE_noblock_obuf_4_2_943_wire;
      req <= phi_stmt_939_req_0 & phi_stmt_939_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_939",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_939_ack_0,
          idata => idata,
          odata => pkt_4_e_word_939,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_939
    phi_stmt_944: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_946_wire_constant & next_active_packet_1027_947_buffered;
      req <= phi_stmt_944_req_0 & phi_stmt_944_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_944",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_944_ack_0,
          idata => idata,
          odata => active_packet_944,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_944
    phi_stmt_948: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_16_950_wire_constant & next_down_counter_1082_951_buffered;
      req <= phi_stmt_948_req_0 & phi_stmt_948_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_948",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_948_ack_0,
          idata => idata,
          odata => down_counter_948,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_948
    phi_stmt_952: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_954_wire_constant & next_pkt_with_priority_1027_955_buffered;
      req <= phi_stmt_952_req_0 & phi_stmt_952_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_952",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_952_ack_0,
          idata => idata,
          odata => pkt_with_priority_952,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_952
    -- flow-through select operator MUX_1001_inst
    MUX_1001_wire <= p2_valid_966 when (EQ_u3_u1_998_wire(0) /=  '0') else konst_1000_wire_constant;
    -- flow-through select operator MUX_1008_inst
    MUX_1008_wire <= p3_valid_971 when (EQ_u3_u1_1005_wire(0) /=  '0') else konst_1007_wire_constant;
    -- flow-through select operator MUX_1014_inst
    MUX_1014_wire <= p4_valid_976 when (EQ_u3_u1_1011_wire(0) /=  '0') else konst_1013_wire_constant;
    -- flow-through select operator MUX_1035_inst
    MUX_1035_wire <= slice_1033_wire when (EQ_u3_u1_1031_wire(0) /=  '0') else konst_1034_wire_constant;
    -- flow-through select operator MUX_1042_inst
    MUX_1042_wire <= slice_1040_wire when (EQ_u3_u1_1038_wire(0) /=  '0') else konst_1041_wire_constant;
    -- flow-through select operator MUX_1050_inst
    MUX_1050_wire <= slice_1048_wire when (EQ_u3_u1_1046_wire(0) /=  '0') else konst_1049_wire_constant;
    -- flow-through select operator MUX_1057_inst
    MUX_1057_wire <= slice_1055_wire when (EQ_u3_u1_1053_wire(0) /=  '0') else konst_1056_wire_constant;
    -- flow-through select operator MUX_1080_inst
    MUX_1080_wire <= SUB_u16_u16_1078_wire when (valid_active_pkt_word_read_1017(0) /=  '0') else down_counter_948;
    -- flow-through select operator MUX_1081_inst
    next_down_counter_1082 <= SUB_u16_u16_1074_wire when (started_new_packet_1069(0) /=  '0') else MUX_1080_wire;
    -- flow-through select operator MUX_1133_inst
    MUX_1133_wire <= slice_1130_wire when (EQ_u3_u1_1128_wire(0) /=  '0') else slice_1132_wire;
    -- flow-through select operator MUX_1134_inst
    MUX_1134_wire <= slice_1125_wire when (EQ_u3_u1_1123_wire(0) /=  '0') else MUX_1133_wire;
    -- flow-through select operator MUX_1135_inst
    data_to_out_1136 <= slice_1120_wire when (EQ_u3_u1_1118_wire(0) /=  '0') else MUX_1134_wire;
    -- flow-through select operator MUX_1143_inst
    MUX_1143_wire <= p1_valid_961 when (EQ_u3_u1_1140_wire(0) /=  '0') else konst_1142_wire_constant;
    -- flow-through select operator MUX_1149_inst
    MUX_1149_wire <= p2_valid_966 when (EQ_u3_u1_1146_wire(0) /=  '0') else konst_1148_wire_constant;
    -- flow-through select operator MUX_1156_inst
    MUX_1156_wire <= p3_valid_971 when (EQ_u3_u1_1153_wire(0) /=  '0') else konst_1155_wire_constant;
    -- flow-through select operator MUX_1162_inst
    MUX_1162_wire <= p4_valid_976 when (EQ_u3_u1_1159_wire(0) /=  '0') else konst_1161_wire_constant;
    -- flow-through select operator MUX_995_inst
    MUX_995_wire <= p1_valid_961 when (EQ_u3_u1_992_wire(0) /=  '0') else konst_994_wire_constant;
    -- flow-through slice operator slice_1033_inst
    slice_1033_wire <= pkt_1_e_word_924(23 downto 8);
    -- flow-through slice operator slice_1040_inst
    slice_1040_wire <= pkt_2_e_word_929(23 downto 8);
    -- flow-through slice operator slice_1048_inst
    slice_1048_wire <= pkt_3_e_word_934(23 downto 8);
    -- flow-through slice operator slice_1055_inst
    slice_1055_wire <= pkt_4_e_word_939(23 downto 8);
    -- flow-through slice operator slice_1120_inst
    slice_1120_wire <= pkt_1_e_word_924(31 downto 0);
    -- flow-through slice operator slice_1125_inst
    slice_1125_wire <= pkt_2_e_word_929(31 downto 0);
    -- flow-through slice operator slice_1130_inst
    slice_1130_wire <= pkt_3_e_word_934(31 downto 0);
    -- flow-through slice operator slice_1132_inst
    slice_1132_wire <= pkt_4_e_word_939(31 downto 0);
    next_active_packet_1027_947_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1027_947_buf_req_0;
      next_active_packet_1027_947_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1027_947_buf_req_1;
      next_active_packet_1027_947_buf_ack_1<= rack(0);
      next_active_packet_1027_947_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1027_947_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1027_947_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1082_951_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1082_951_buf_req_0;
      next_down_counter_1082_951_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1082_951_buf_req_1;
      next_down_counter_1082_951_buf_ack_1<= rack(0);
      next_down_counter_1082_951_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1082_951_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1082,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1082_951_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_with_priority_1027_955_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_with_priority_1027_955_buf_req_0;
      next_pkt_with_priority_1027_955_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_with_priority_1027_955_buf_req_1;
      next_pkt_with_priority_1027_955_buf_ack_1<= rack(0);
      next_pkt_with_priority_1027_955_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_with_priority_1027_955_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_with_priority_1027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_with_priority_1027_955_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_922_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1180_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_922_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_922_branch_req_0,
          ack0 => do_while_stmt_922_branch_ack_0,
          ack1 => do_while_stmt_922_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1068_inst
    process(NEQ_u3_u1_1064_wire, EQ_u16_u1_1067_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u3_u1_1064_wire, EQ_u16_u1_1067_wire, tmp_var);
      started_new_packet_1069 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_960_inst
    process(pkt_1_e_word_924) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_924, konst_959_wire_constant, tmp_var);
      p1_valid_961 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_965_inst
    process(pkt_2_e_word_929) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_929, konst_964_wire_constant, tmp_var);
      p2_valid_966 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_970_inst
    process(pkt_3_e_word_934) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_934, konst_969_wire_constant, tmp_var);
      p3_valid_971 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_975_inst
    process(pkt_4_e_word_939) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_939, konst_974_wire_constant, tmp_var);
      p4_valid_976 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1067_inst
    process(down_counter_948) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_948, konst_1066_wire_constant, tmp_var);
      EQ_u16_u1_1067_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1005_inst
    process(active_packet_944) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_944, konst_1004_wire_constant, tmp_var);
      EQ_u3_u1_1005_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1011_inst
    process(active_packet_944) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_944, konst_1010_wire_constant, tmp_var);
      EQ_u3_u1_1011_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1031_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1030_wire_constant, tmp_var);
      EQ_u3_u1_1031_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1038_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1037_wire_constant, tmp_var);
      EQ_u3_u1_1038_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1046_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1045_wire_constant, tmp_var);
      EQ_u3_u1_1046_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1053_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1052_wire_constant, tmp_var);
      EQ_u3_u1_1053_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1088_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1087_wire_constant, tmp_var);
      EQ_u3_u1_1088_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1096_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1095_wire_constant, tmp_var);
      EQ_u3_u1_1096_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1104_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1103_wire_constant, tmp_var);
      EQ_u3_u1_1104_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1112_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1111_wire_constant, tmp_var);
      EQ_u3_u1_1112_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1118_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1117_wire_constant, tmp_var);
      EQ_u3_u1_1118_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1123_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1122_wire_constant, tmp_var);
      EQ_u3_u1_1123_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1128_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1127_wire_constant, tmp_var);
      EQ_u3_u1_1128_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1140_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1139_wire_constant, tmp_var);
      EQ_u3_u1_1140_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1146_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1145_wire_constant, tmp_var);
      EQ_u3_u1_1146_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1153_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1152_wire_constant, tmp_var);
      EQ_u3_u1_1153_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1159_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1027, konst_1158_wire_constant, tmp_var);
      EQ_u3_u1_1159_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_992_inst
    process(active_packet_944) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_944, konst_991_wire_constant, tmp_var);
      EQ_u3_u1_992_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_998_inst
    process(active_packet_944) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_944, konst_997_wire_constant, tmp_var);
      EQ_u3_u1_998_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_1064_inst
    process(next_active_packet_1027) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_1027, konst_1063_wire_constant, tmp_var);
      NEQ_u3_u1_1064_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1085_inst
    process(p1_valid_961) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_961, tmp_var);
      NOT_u1_u1_1085_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1093_inst
    process(p2_valid_966) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_966, tmp_var);
      NOT_u1_u1_1093_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1101_inst
    process(p3_valid_971) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_971, tmp_var);
      NOT_u1_u1_1101_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1109_inst
    process(p4_valid_976) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_976, tmp_var);
      NOT_u1_u1_1109_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_1043_inst
    process(MUX_1035_wire, MUX_1042_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1035_wire, MUX_1042_wire, tmp_var);
      OR_u16_u16_1043_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1058_inst
    process(MUX_1050_wire, MUX_1057_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1050_wire, MUX_1057_wire, tmp_var);
      OR_u16_u16_1058_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1059_inst
    process(OR_u16_u16_1043_wire, OR_u16_u16_1058_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u16_u16_1043_wire, OR_u16_u16_1058_wire, tmp_var);
      valid_active_pkt_length_1060 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1002_inst
    process(MUX_995_wire, MUX_1001_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_995_wire, MUX_1001_wire, tmp_var);
      OR_u1_u1_1002_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1015_inst
    process(MUX_1008_wire, MUX_1014_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1008_wire, MUX_1014_wire, tmp_var);
      OR_u1_u1_1015_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1016_inst
    process(OR_u1_u1_1002_wire, OR_u1_u1_1015_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1002_wire, OR_u1_u1_1015_wire, tmp_var);
      valid_active_pkt_word_read_1017 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1089_inst
    process(NOT_u1_u1_1085_wire, EQ_u3_u1_1088_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1085_wire, EQ_u3_u1_1088_wire, tmp_var);
      read_from_1_1090 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1097_inst
    process(NOT_u1_u1_1093_wire, EQ_u3_u1_1096_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1093_wire, EQ_u3_u1_1096_wire, tmp_var);
      read_from_2_1098 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1105_inst
    process(NOT_u1_u1_1101_wire, EQ_u3_u1_1104_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1101_wire, EQ_u3_u1_1104_wire, tmp_var);
      read_from_3_1106 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1113_inst
    process(NOT_u1_u1_1109_wire, EQ_u3_u1_1112_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1109_wire, EQ_u3_u1_1112_wire, tmp_var);
      read_from_4_1114 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1150_inst
    process(MUX_1143_wire, MUX_1149_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1143_wire, MUX_1149_wire, tmp_var);
      OR_u1_u1_1150_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1163_inst
    process(MUX_1156_wire, MUX_1162_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1156_wire, MUX_1162_wire, tmp_var);
      OR_u1_u1_1163_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1164_inst
    process(OR_u1_u1_1150_wire, OR_u1_u1_1163_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1150_wire, OR_u1_u1_1163_wire, tmp_var);
      send_flag_1165 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1074_inst
    process(valid_active_pkt_length_1060) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(valid_active_pkt_length_1060, konst_1073_wire_constant, tmp_var);
      SUB_u16_u16_1074_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1078_inst
    process(down_counter_948) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_948, konst_1077_wire_constant, tmp_var);
      SUB_u16_u16_1078_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_2_928_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_2_928_inst_req_0;
      RPIPE_noblock_obuf_1_2_928_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_2_928_inst_req_1;
      RPIPE_noblock_obuf_1_2_928_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1090(0);
      RPIPE_noblock_obuf_1_2_928_wire <= data_out(32 downto 0);
      noblock_obuf_1_2_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_2_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_2_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_2_pipe_read_req(0),
          oack => noblock_obuf_1_2_pipe_read_ack(0),
          odata => noblock_obuf_1_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_2_933_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_2_933_inst_req_0;
      RPIPE_noblock_obuf_2_2_933_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_2_933_inst_req_1;
      RPIPE_noblock_obuf_2_2_933_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1098(0);
      RPIPE_noblock_obuf_2_2_933_wire <= data_out(32 downto 0);
      noblock_obuf_2_2_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_2_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_2_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_2_pipe_read_req(0),
          oack => noblock_obuf_2_2_pipe_read_ack(0),
          odata => noblock_obuf_2_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_2_938_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_2_938_inst_req_0;
      RPIPE_noblock_obuf_3_2_938_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_2_938_inst_req_1;
      RPIPE_noblock_obuf_3_2_938_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1106(0);
      RPIPE_noblock_obuf_3_2_938_wire <= data_out(32 downto 0);
      noblock_obuf_3_2_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_2_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_2_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_2_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_2_pipe_read_req(0),
          oack => noblock_obuf_3_2_pipe_read_ack(0),
          odata => noblock_obuf_3_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_2_943_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_2_943_inst_req_0;
      RPIPE_noblock_obuf_4_2_943_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_2_943_inst_req_1;
      RPIPE_noblock_obuf_4_2_943_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1114(0);
      RPIPE_noblock_obuf_4_2_943_wire <= data_out(32 downto 0);
      noblock_obuf_4_2_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_2_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_2_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_2_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_2_pipe_read_req(0),
          oack => noblock_obuf_4_2_pipe_read_ack(0),
          odata => noblock_obuf_4_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_2_1167_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_2_1167_inst_req_0;
      WPIPE_out_data_2_1167_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_2_1167_inst_req_1;
      WPIPE_out_data_2_1167_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1165(0);
      data_in <= data_to_out_1136;
      out_data_2_write_0_gI: SplitGuardInterface generic map(name => "out_data_2_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_2_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_2", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_2_pipe_write_req(0),
          oack => out_data_2_pipe_write_ack(0),
          odata => out_data_2_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_2524: prioritySelect_Volatile port map(down_counter => down_counter_948, active_packet => active_packet_944, pkt_with_priority => pkt_with_priority_952, p1_valid => p1_valid_961, p2_valid => p2_valid_966, p3_valid => p3_valid_971, p4_valid => p4_valid_976, next_active_packet => next_active_packet_1027, next_pkt_with_priority => next_pkt_with_priority_1027); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_2_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_3_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_3_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_3_Daemon;
architecture outputPort_3_Daemon_arch of outputPort_3_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_3_Daemon_CP_1538_start: Boolean;
  signal outputPort_3_Daemon_CP_1538_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(15 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_with_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_with_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal WPIPE_out_data_3_1430_inst_req_1 : boolean;
  signal next_pkt_with_priority_1290_1218_buf_ack_1 : boolean;
  signal phi_stmt_1211_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_3_1206_inst_ack_1 : boolean;
  signal next_active_packet_1290_1210_buf_req_0 : boolean;
  signal phi_stmt_1207_req_1 : boolean;
  signal phi_stmt_1211_ack_0 : boolean;
  signal phi_stmt_1207_ack_0 : boolean;
  signal WPIPE_out_data_3_1430_inst_ack_0 : boolean;
  signal phi_stmt_1211_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_3_1206_inst_req_0 : boolean;
  signal next_active_packet_1290_1210_buf_ack_0 : boolean;
  signal next_pkt_with_priority_1290_1218_buf_req_1 : boolean;
  signal next_pkt_with_priority_1290_1218_buf_req_0 : boolean;
  signal WPIPE_out_data_3_1430_inst_ack_1 : boolean;
  signal WPIPE_out_data_3_1430_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_3_1206_inst_ack_0 : boolean;
  signal do_while_stmt_1185_branch_ack_0 : boolean;
  signal next_pkt_with_priority_1290_1218_buf_ack_0 : boolean;
  signal phi_stmt_1207_req_0 : boolean;
  signal next_down_counter_1345_1214_buf_req_0 : boolean;
  signal next_down_counter_1345_1214_buf_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_3_1206_inst_req_1 : boolean;
  signal next_active_packet_1290_1210_buf_req_1 : boolean;
  signal do_while_stmt_1185_branch_ack_1 : boolean;
  signal next_down_counter_1345_1214_buf_req_1 : boolean;
  signal next_down_counter_1345_1214_buf_ack_1 : boolean;
  signal next_active_packet_1290_1210_buf_ack_1 : boolean;
  signal phi_stmt_1215_req_1 : boolean;
  signal phi_stmt_1215_req_0 : boolean;
  signal phi_stmt_1215_ack_0 : boolean;
  signal do_while_stmt_1185_branch_req_0 : boolean;
  signal phi_stmt_1187_req_1 : boolean;
  signal phi_stmt_1187_req_0 : boolean;
  signal phi_stmt_1187_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1191_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1191_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1191_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_3_1191_inst_ack_1 : boolean;
  signal phi_stmt_1192_req_1 : boolean;
  signal phi_stmt_1192_req_0 : boolean;
  signal phi_stmt_1192_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1196_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1196_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1196_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_3_1196_inst_ack_1 : boolean;
  signal phi_stmt_1197_req_1 : boolean;
  signal phi_stmt_1197_req_0 : boolean;
  signal phi_stmt_1197_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_3_1201_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_3_1201_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_3_1201_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_3_1201_inst_ack_1 : boolean;
  signal phi_stmt_1202_req_1 : boolean;
  signal phi_stmt_1202_req_0 : boolean;
  signal phi_stmt_1202_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_3_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_3_Daemon_CP_1538_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_3_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_3_Daemon_CP_1538: Block -- control-path 
    signal outputPort_3_Daemon_CP_1538_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_3_Daemon_CP_1538_elements(0) <= outputPort_3_Daemon_CP_1538_start;
    outputPort_3_Daemon_CP_1538_symbol <= outputPort_3_Daemon_CP_1538_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1184/$entry
      -- CP-element group 0: 	 branch_block_stmt_1184/branch_block_stmt_1184__entry__
      -- CP-element group 0: 	 branch_block_stmt_1184/do_while_stmt_1185__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1184/$exit
      -- CP-element group 1: 	 branch_block_stmt_1184/branch_block_stmt_1184__exit__
      -- CP-element group 1: 	 branch_block_stmt_1184/do_while_stmt_1185__exit__
      -- 
    outputPort_3_Daemon_CP_1538_elements(1) <= outputPort_3_Daemon_CP_1538_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1184/do_while_stmt_1185/$entry
      -- CP-element group 2: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185__entry__
      -- 
    outputPort_3_Daemon_CP_1538_elements(2) <= outputPort_3_Daemon_CP_1538_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185__exit__
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1184/do_while_stmt_1185/loop_back
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	159 
    -- CP-element group 5: 	160 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1184/do_while_stmt_1185/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1184/do_while_stmt_1185/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1184/do_while_stmt_1185/condition_done
      -- 
    outputPort_3_Daemon_CP_1538_elements(5) <= outputPort_3_Daemon_CP_1538_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1184/do_while_stmt_1185/loop_body_done
      -- 
    outputPort_3_Daemon_CP_1538_elements(6) <= outputPort_3_Daemon_CP_1538_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	61 
    -- CP-element group 7: 	82 
    -- CP-element group 7: 	103 
    -- CP-element group 7: 	122 
    -- CP-element group 7: 	141 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/back_edge_to_loop_body
      -- 
    outputPort_3_Daemon_CP_1538_elements(7) <= outputPort_3_Daemon_CP_1538_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	63 
    -- CP-element group 8: 	84 
    -- CP-element group 8: 	105 
    -- CP-element group 8: 	124 
    -- CP-element group 8: 	143 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/first_time_through_loop_body
      -- 
    outputPort_3_Daemon_CP_1538_elements(8) <= outputPort_3_Daemon_CP_1538_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	76 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	97 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	116 
    -- CP-element group 9: 	117 
    -- CP-element group 9: 	135 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	157 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/loop_body_start
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	157 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/condition_evaluated
      -- 
    condition_evaluated_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(10), ack => do_while_stmt_1185_branch_req_0); -- 
    outputPort_3_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(14) & outputPort_3_Daemon_CP_1538_elements(157);
      gj_outputPort_3_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	97 
    -- CP-element group 11: 	116 
    -- CP-element group 11: 	135 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11: 	99 
    -- CP-element group 11: 	118 
    -- CP-element group 11: 	137 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_sample_start__ps
      -- 
    outputPort_3_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(15) & outputPort_3_Daemon_CP_1538_elements(34) & outputPort_3_Daemon_CP_1538_elements(55) & outputPort_3_Daemon_CP_1538_elements(76) & outputPort_3_Daemon_CP_1538_elements(97) & outputPort_3_Daemon_CP_1538_elements(116) & outputPort_3_Daemon_CP_1538_elements(135) & outputPort_3_Daemon_CP_1538_elements(14);
      gj_outputPort_3_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	58 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	100 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	138 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	55 
    -- CP-element group 12: 	76 
    -- CP-element group 12: 	97 
    -- CP-element group 12: 	116 
    -- CP-element group 12: 	135 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_sample_completed_
      -- 
    outputPort_3_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(17) & outputPort_3_Daemon_CP_1538_elements(37) & outputPort_3_Daemon_CP_1538_elements(58) & outputPort_3_Daemon_CP_1538_elements(79) & outputPort_3_Daemon_CP_1538_elements(100) & outputPort_3_Daemon_CP_1538_elements(119) & outputPort_3_Daemon_CP_1538_elements(138);
      gj_outputPort_3_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	77 
    -- CP-element group 13: 	98 
    -- CP-element group 13: 	117 
    -- CP-element group 13: 	136 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	59 
    -- CP-element group 13: 	80 
    -- CP-element group 13: 	101 
    -- CP-element group 13: 	120 
    -- CP-element group 13: 	139 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_update_start__ps
      -- 
    outputPort_3_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(16) & outputPort_3_Daemon_CP_1538_elements(35) & outputPort_3_Daemon_CP_1538_elements(56) & outputPort_3_Daemon_CP_1538_elements(77) & outputPort_3_Daemon_CP_1538_elements(98) & outputPort_3_Daemon_CP_1538_elements(117) & outputPort_3_Daemon_CP_1538_elements(136);
      gj_outputPort_3_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	102 
    -- CP-element group 14: 	121 
    -- CP-element group 14: 	140 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_3_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(18) & outputPort_3_Daemon_CP_1538_elements(39) & outputPort_3_Daemon_CP_1538_elements(60) & outputPort_3_Daemon_CP_1538_elements(81) & outputPort_3_Daemon_CP_1538_elements(102) & outputPort_3_Daemon_CP_1538_elements(121) & outputPort_3_Daemon_CP_1538_elements(140);
      gj_outputPort_3_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	154 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(19) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_loopback_sample_req_ps
      -- 
    phi_stmt_1187_loopback_sample_req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1187_loopback_sample_req_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(20), ack => phi_stmt_1187_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(21) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_entry_sample_req_ps
      -- 
    phi_stmt_1187_entry_sample_req_1580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1187_entry_sample_req_1580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(22), ack => phi_stmt_1187_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1187_phi_mux_ack_ps
      -- 
    phi_stmt_1187_phi_mux_ack_1583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1187_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1189_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1189_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1189_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1189_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1189_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1189_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1189_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(26) <= outputPort_3_Daemon_CP_1538_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1189_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(25), ack => outputPort_3_Daemon_CP_1538_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	33 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_Sample/rr
      -- 
    rr_1604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(30), ack => RPIPE_noblock_obuf_1_3_1191_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(28) & outputPort_3_Daemon_CP_1538_elements(33);
      gj_outputPort_3_Daemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: 	32 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_Update/cr
      -- 
    cr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(31), ack => RPIPE_noblock_obuf_1_3_1191_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(29) & outputPort_3_Daemon_CP_1538_elements(32);
      gj_outputPort_3_Daemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	31 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_Sample/ra
      -- 
    ra_1605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_3_1191_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	30 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_1_3_1191_Update/ca
      -- 
    ca_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_3_1191_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	155 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(36) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(38) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: 	154 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(40) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_loopback_sample_req_ps
      -- 
    phi_stmt_1192_loopback_sample_req_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1192_loopback_sample_req_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(41), ack => phi_stmt_1192_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(42) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_entry_sample_req_ps
      -- 
    phi_stmt_1192_entry_sample_req_1624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1192_entry_sample_req_1624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(43), ack => phi_stmt_1192_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1192_phi_mux_ack_ps
      -- 
    phi_stmt_1192_phi_mux_ack_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1192_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1194_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1194_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1194_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1194_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1194_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1194_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1194_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(47) <= outputPort_3_Daemon_CP_1538_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1194_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(46), ack => outputPort_3_Daemon_CP_1538_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_Sample/rr
      -- 
    rr_1648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(51), ack => RPIPE_noblock_obuf_2_3_1196_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(49) & outputPort_3_Daemon_CP_1538_elements(54);
      gj_outputPort_3_Daemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	53 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_Update/cr
      -- 
    cr_1653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(52), ack => RPIPE_noblock_obuf_2_3_1196_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(50) & outputPort_3_Daemon_CP_1538_elements(53);
      gj_outputPort_3_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	52 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_Sample/ra
      -- 
    ra_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_3_1196_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_2_3_1196_Update/ca
      -- 
    ca_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_3_1196_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	155 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(57) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(59) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	14 
    -- CP-element group 60: 	154 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(61) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_loopback_sample_req_ps
      -- 
    phi_stmt_1197_loopback_sample_req_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1197_loopback_sample_req_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(62), ack => phi_stmt_1197_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(63) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_entry_sample_req_ps
      -- 
    phi_stmt_1197_entry_sample_req_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1197_entry_sample_req_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(64), ack => phi_stmt_1197_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1197_phi_mux_ack_ps
      -- 
    phi_stmt_1197_phi_mux_ack_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1197_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1199_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1199_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1199_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1199_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1199_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1199_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1199_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(68) <= outputPort_3_Daemon_CP_1538_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1199_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(67), ack => outputPort_3_Daemon_CP_1538_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	75 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_Sample/rr
      -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(72), ack => RPIPE_noblock_obuf_3_3_1201_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(70) & outputPort_3_Daemon_CP_1538_elements(75);
      gj_outputPort_3_Daemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	74 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_update_start_
      -- CP-element group 73: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_Update/cr
      -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(73), ack => RPIPE_noblock_obuf_3_3_1201_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(71) & outputPort_3_Daemon_CP_1538_elements(74);
      gj_outputPort_3_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	73 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_Sample/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_3_1201_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	72 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_3_3_1201_Update/ca
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_3_1201_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	9 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	12 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	11 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	155 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	11 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(78) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	12 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	13 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(80) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: 	154 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	7 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(82) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_loopback_sample_req_ps
      -- 
    phi_stmt_1202_loopback_sample_req_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1202_loopback_sample_req_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(83), ack => phi_stmt_1202_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(84) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_entry_sample_req_ps
      -- 
    phi_stmt_1202_entry_sample_req_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1202_entry_sample_req_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(85), ack => phi_stmt_1202_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_phi_mux_ack_ps
      -- CP-element group 86: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1202_phi_mux_ack
      -- 
    phi_stmt_1202_phi_mux_ack_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1202_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1204_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1204_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1204_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1204_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1204_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1204_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1204_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(89) <= outputPort_3_Daemon_CP_1538_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_33_1204_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(88), ack => outputPort_3_Daemon_CP_1538_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	96 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_Sample/$entry
      -- 
    rr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(93), ack => RPIPE_noblock_obuf_4_3_1206_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(91) & outputPort_3_Daemon_CP_1538_elements(96);
      gj_outputPort_3_Daemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	95 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_Update/cr
      -- 
    cr_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(94), ack => RPIPE_noblock_obuf_4_3_1206_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(92) & outputPort_3_Daemon_CP_1538_elements(95);
      gj_outputPort_3_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	94 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_sample_completed__ps
      -- 
    ra_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_3_1206_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	93 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/RPIPE_noblock_obuf_4_3_1206_update_completed__ps
      -- 
    ca_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_3_1206_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	9 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	11 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	155 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	13 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	11 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(99) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	12 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	13 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(101) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	14 
    -- CP-element group 102: 	154 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_update_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	7 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(103) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_loopback_sample_req
      -- CP-element group 104: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_loopback_sample_req_ps
      -- 
    phi_stmt_1207_loopback_sample_req_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1207_loopback_sample_req_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(104), ack => phi_stmt_1207_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	8 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(105) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_entry_sample_req_ps
      -- CP-element group 106: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_entry_sample_req
      -- 
    phi_stmt_1207_entry_sample_req_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1207_entry_sample_req_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(106), ack => phi_stmt_1207_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1207_phi_mux_ack_ps
      -- 
    phi_stmt_1207_phi_mux_ack_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1207_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_3_1209_sample_start__ps
      -- CP-element group 108: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_3_1209_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_3_1209_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_3_1209_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_3_1209_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_3_1209_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_3_1209_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(110) <= outputPort_3_Daemon_CP_1538_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_3_1209_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(109), ack => outputPort_3_Daemon_CP_1538_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_Sample/req
      -- CP-element group 112: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_sample_start__ps
      -- CP-element group 112: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_sample_start_
      -- 
    req_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(112), ack => next_active_packet_1290_1210_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_Update/req
      -- CP-element group 113: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_update_start__ps
      -- 
    req_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(113), ack => next_active_packet_1290_1210_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_sample_completed_
      -- 
    ack_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1290_1210_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(114)); -- 
    -- CP-element group 115:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_Update/ack
      -- CP-element group 115: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_active_packet_1210_update_completed__ps
      -- 
    ack_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1290_1210_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(115)); -- 
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	9 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	12 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	11 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	9 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	155 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	13 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	11 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(118) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	12 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	13 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(120) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	14 
    -- CP-element group 121: 	154 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	7 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(122) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_loopback_sample_req
      -- CP-element group 123: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_loopback_sample_req_ps
      -- 
    phi_stmt_1211_loopback_sample_req_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1211_loopback_sample_req_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(123), ack => phi_stmt_1211_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(124) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_entry_sample_req
      -- CP-element group 125: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_entry_sample_req_ps
      -- 
    phi_stmt_1211_entry_sample_req_1800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1211_entry_sample_req_1800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(125), ack => phi_stmt_1211_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_phi_mux_ack
      -- CP-element group 126: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1211_phi_mux_ack_ps
      -- 
    phi_stmt_1211_phi_mux_ack_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1211_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_16_1213_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_16_1213_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_16_1213_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_16_1213_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_16_1213_update_start_
      -- CP-element group 128: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_16_1213_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_16_1213_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(129) <= outputPort_3_Daemon_CP_1538_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_ZERO_16_1213_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(128), ack => outputPort_3_Daemon_CP_1538_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_sample_start__ps
      -- CP-element group 131: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_Sample/req
      -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(131), ack => next_down_counter_1345_1214_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_update_start__ps
      -- CP-element group 132: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_update_start_
      -- CP-element group 132: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_Update/req
      -- 
    req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(132), ack => next_down_counter_1345_1214_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_Sample/ack
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1345_1214_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(133)); -- 
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_down_counter_1214_Update/ack
      -- 
    ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1345_1214_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	9 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	11 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	155 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	13 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(137) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	12 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	13 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(139) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	14 
    -- CP-element group 140: 	154 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(141) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_loopback_sample_req_ps
      -- 
    phi_stmt_1215_loopback_sample_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1215_loopback_sample_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(142), ack => phi_stmt_1215_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(143) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_entry_sample_req_ps
      -- 
    phi_stmt_1215_entry_sample_req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1215_entry_sample_req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(144), ack => phi_stmt_1215_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/phi_stmt_1215_phi_mux_ack_ps
      -- 
    phi_stmt_1215_phi_mux_ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1215_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/konst_1217_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/konst_1217_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/konst_1217_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/konst_1217_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/konst_1217_update_start_
      -- CP-element group 147: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/konst_1217_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/konst_1217_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(148) <= outputPort_3_Daemon_CP_1538_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/konst_1217_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(147), ack => outputPort_3_Daemon_CP_1538_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_sample_start_
      -- 
    req_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(150), ack => next_pkt_with_priority_1290_1218_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_Update/req
      -- 
    req_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(151), ack => next_pkt_with_priority_1290_1218_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_Sample/ack
      -- 
    ack_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_with_priority_1290_1218_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/R_next_pkt_with_priority_1218_update_completed_
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_with_priority_1290_1218_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	18 
    -- CP-element group 154: 	39 
    -- CP-element group 154: 	60 
    -- CP-element group 154: 	81 
    -- CP-element group 154: 	102 
    -- CP-element group 154: 	121 
    -- CP-element group 154: 	140 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_Sample/req
      -- CP-element group 154: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_sample_start_
      -- 
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(154), ack => WPIPE_out_data_3_1430_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(18) & outputPort_3_Daemon_CP_1538_elements(39) & outputPort_3_Daemon_CP_1538_elements(60) & outputPort_3_Daemon_CP_1538_elements(81) & outputPort_3_Daemon_CP_1538_elements(102) & outputPort_3_Daemon_CP_1538_elements(121) & outputPort_3_Daemon_CP_1538_elements(140) & outputPort_3_Daemon_CP_1538_elements(156);
      gj_outputPort_3_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	35 
    -- CP-element group 155: 	56 
    -- CP-element group 155: 	77 
    -- CP-element group 155: 	98 
    -- CP-element group 155: 	117 
    -- CP-element group 155: 	136 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_Update/req
      -- CP-element group 155: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_update_start_
      -- 
    ack_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3_1430_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(155)); -- 
    req_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(155), ack => WPIPE_out_data_3_1430_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_Update/ack
      -- CP-element group 156: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/WPIPE_out_data_3_1430_update_completed_
      -- 
    ack_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3_1430_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(9), ack => outputPort_3_Daemon_CP_1538_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	12 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1184/do_while_stmt_1185/do_while_stmt_1185_loop_body/$exit
      -- 
    outputPort_3_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(12) & outputPort_3_Daemon_CP_1538_elements(156);
      gj_outputPort_3_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_1184/do_while_stmt_1185/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_1184/do_while_stmt_1185/loop_exit/ack
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1185_branch_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1184/do_while_stmt_1185/loop_taken/$exit
      -- CP-element group 160: 	 branch_block_stmt_1184/do_while_stmt_1185/loop_taken/ack
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1185_branch_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1184/do_while_stmt_1185/$exit
      -- 
    outputPort_3_Daemon_CP_1538_elements(161) <= outputPort_3_Daemon_CP_1538_elements(3);
    outputPort_3_Daemon_do_while_stmt_1185_terminator_1899: loop_terminator -- 
      generic map (name => " outputPort_3_Daemon_do_while_stmt_1185_terminator_1899", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_3_Daemon_CP_1538_elements(6),loop_continue => outputPort_3_Daemon_CP_1538_elements(160),loop_terminate => outputPort_3_Daemon_CP_1538_elements(159),loop_back => outputPort_3_Daemon_CP_1538_elements(4),loop_exit => outputPort_3_Daemon_CP_1538_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1187_phi_seq_1611_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(21);
      outputPort_3_Daemon_CP_1538_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(24);
      outputPort_3_Daemon_CP_1538_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(26);
      outputPort_3_Daemon_CP_1538_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(19);
      outputPort_3_Daemon_CP_1538_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(32);
      outputPort_3_Daemon_CP_1538_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(33);
      outputPort_3_Daemon_CP_1538_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1187_phi_seq_1611 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1187_phi_seq_1611") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(11), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(17), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(13), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(18), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1192_phi_seq_1655_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(42);
      outputPort_3_Daemon_CP_1538_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(45);
      outputPort_3_Daemon_CP_1538_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(47);
      outputPort_3_Daemon_CP_1538_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(40);
      outputPort_3_Daemon_CP_1538_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(53);
      outputPort_3_Daemon_CP_1538_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(54);
      outputPort_3_Daemon_CP_1538_elements(41) <= phi_mux_reqs(1);
      phi_stmt_1192_phi_seq_1655 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1192_phi_seq_1655") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(36), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(37), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(38), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(39), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1197_phi_seq_1699_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(63);
      outputPort_3_Daemon_CP_1538_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(66);
      outputPort_3_Daemon_CP_1538_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(68);
      outputPort_3_Daemon_CP_1538_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(61);
      outputPort_3_Daemon_CP_1538_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(74);
      outputPort_3_Daemon_CP_1538_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(75);
      outputPort_3_Daemon_CP_1538_elements(62) <= phi_mux_reqs(1);
      phi_stmt_1197_phi_seq_1699 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1197_phi_seq_1699") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(57), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(58), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(59), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(60), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1202_phi_seq_1743_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(84);
      outputPort_3_Daemon_CP_1538_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(87);
      outputPort_3_Daemon_CP_1538_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(89);
      outputPort_3_Daemon_CP_1538_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(82);
      outputPort_3_Daemon_CP_1538_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(95);
      outputPort_3_Daemon_CP_1538_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(96);
      outputPort_3_Daemon_CP_1538_elements(83) <= phi_mux_reqs(1);
      phi_stmt_1202_phi_seq_1743 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1202_phi_seq_1743") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(78), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(79), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(80), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(81), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1207_phi_seq_1787_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(105);
      outputPort_3_Daemon_CP_1538_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(108);
      outputPort_3_Daemon_CP_1538_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(110);
      outputPort_3_Daemon_CP_1538_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(103);
      outputPort_3_Daemon_CP_1538_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(114);
      outputPort_3_Daemon_CP_1538_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(115);
      outputPort_3_Daemon_CP_1538_elements(104) <= phi_mux_reqs(1);
      phi_stmt_1207_phi_seq_1787 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1207_phi_seq_1787") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(99), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(100), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(101), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(102), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1211_phi_seq_1831_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(124);
      outputPort_3_Daemon_CP_1538_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(127);
      outputPort_3_Daemon_CP_1538_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(129);
      outputPort_3_Daemon_CP_1538_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(122);
      outputPort_3_Daemon_CP_1538_elements(131)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(133);
      outputPort_3_Daemon_CP_1538_elements(132)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(134);
      outputPort_3_Daemon_CP_1538_elements(123) <= phi_mux_reqs(1);
      phi_stmt_1211_phi_seq_1831 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1211_phi_seq_1831") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(118), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(119), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(120), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(121), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1215_phi_seq_1875_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(143);
      outputPort_3_Daemon_CP_1538_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(146);
      outputPort_3_Daemon_CP_1538_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(148);
      outputPort_3_Daemon_CP_1538_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(141);
      outputPort_3_Daemon_CP_1538_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(152);
      outputPort_3_Daemon_CP_1538_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(153);
      outputPort_3_Daemon_CP_1538_elements(142) <= phi_mux_reqs(1);
      phi_stmt_1215_phi_seq_1875 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1215_phi_seq_1875") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(137), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(138), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(139), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(140), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1563_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_3_Daemon_CP_1538_elements(7);
        preds(1)  <= outputPort_3_Daemon_CP_1538_elements(8);
        entry_tmerge_1563 : transition_merge -- 
          generic map(name => " entry_tmerge_1563")
          port map (preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u16_u1_1330_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1255_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1261_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1268_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1274_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1294_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1301_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1309_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1316_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1351_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1359_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1367_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1375_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1381_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1386_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1391_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1403_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1409_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1416_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1422_wire : std_logic_vector(0 downto 0);
    signal MUX_1258_wire : std_logic_vector(0 downto 0);
    signal MUX_1264_wire : std_logic_vector(0 downto 0);
    signal MUX_1271_wire : std_logic_vector(0 downto 0);
    signal MUX_1277_wire : std_logic_vector(0 downto 0);
    signal MUX_1298_wire : std_logic_vector(15 downto 0);
    signal MUX_1305_wire : std_logic_vector(15 downto 0);
    signal MUX_1313_wire : std_logic_vector(15 downto 0);
    signal MUX_1320_wire : std_logic_vector(15 downto 0);
    signal MUX_1343_wire : std_logic_vector(15 downto 0);
    signal MUX_1396_wire : std_logic_vector(31 downto 0);
    signal MUX_1397_wire : std_logic_vector(31 downto 0);
    signal MUX_1406_wire : std_logic_vector(0 downto 0);
    signal MUX_1412_wire : std_logic_vector(0 downto 0);
    signal MUX_1419_wire : std_logic_vector(0 downto 0);
    signal MUX_1425_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_1327_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1348_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1356_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1364_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1372_wire : std_logic_vector(0 downto 0);
    signal OR_u16_u16_1306_wire : std_logic_vector(15 downto 0);
    signal OR_u16_u16_1321_wire : std_logic_vector(15 downto 0);
    signal OR_u1_u1_1265_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1278_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1413_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1426_wire : std_logic_vector(0 downto 0);
    signal RPIPE_noblock_obuf_1_3_1191_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_3_1196_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_3_1201_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_3_1206_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_16_1213_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_33_1189_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1194_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1199_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1204_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1209_wire_constant : std_logic_vector(2 downto 0);
    signal SUB_u16_u16_1337_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_1341_wire : std_logic_vector(15 downto 0);
    signal active_packet_1207 : std_logic_vector(2 downto 0);
    signal data_to_out_1399 : std_logic_vector(31 downto 0);
    signal down_counter_1211 : std_logic_vector(15 downto 0);
    signal konst_1217_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1222_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1227_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1232_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1237_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1254_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1257_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1260_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1263_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1267_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1270_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1273_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1276_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1293_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1297_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1300_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1304_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1308_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1312_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1315_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1319_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1326_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1329_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1336_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1340_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1350_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1358_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1366_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1374_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1380_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1385_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1390_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1402_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1405_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1408_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1411_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1415_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1418_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1421_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1424_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1443_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1290 : std_logic_vector(2 downto 0);
    signal next_active_packet_1290_1210_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_1345 : std_logic_vector(15 downto 0);
    signal next_down_counter_1345_1214_buffered : std_logic_vector(15 downto 0);
    signal next_pkt_with_priority_1290 : std_logic_vector(2 downto 0);
    signal next_pkt_with_priority_1290_1218_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_1224 : std_logic_vector(0 downto 0);
    signal p2_valid_1229 : std_logic_vector(0 downto 0);
    signal p3_valid_1234 : std_logic_vector(0 downto 0);
    signal p4_valid_1239 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1187 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1192 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1197 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1202 : std_logic_vector(32 downto 0);
    signal pkt_with_priority_1215 : std_logic_vector(2 downto 0);
    signal read_from_1_1353 : std_logic_vector(0 downto 0);
    signal read_from_2_1361 : std_logic_vector(0 downto 0);
    signal read_from_3_1369 : std_logic_vector(0 downto 0);
    signal read_from_4_1377 : std_logic_vector(0 downto 0);
    signal send_flag_1428 : std_logic_vector(0 downto 0);
    signal slice_1296_wire : std_logic_vector(15 downto 0);
    signal slice_1303_wire : std_logic_vector(15 downto 0);
    signal slice_1311_wire : std_logic_vector(15 downto 0);
    signal slice_1318_wire : std_logic_vector(15 downto 0);
    signal slice_1383_wire : std_logic_vector(31 downto 0);
    signal slice_1388_wire : std_logic_vector(31 downto 0);
    signal slice_1393_wire : std_logic_vector(31 downto 0);
    signal slice_1395_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1332 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_length_1323 : std_logic_vector(15 downto 0);
    signal valid_active_pkt_word_read_1280 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_16_1213_wire_constant <= "0000000000000000";
    R_ZERO_33_1189_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1194_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1199_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1204_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1209_wire_constant <= "000";
    konst_1217_wire_constant <= "001";
    konst_1222_wire_constant <= "000000000000000000000000000100000";
    konst_1227_wire_constant <= "000000000000000000000000000100000";
    konst_1232_wire_constant <= "000000000000000000000000000100000";
    konst_1237_wire_constant <= "000000000000000000000000000100000";
    konst_1254_wire_constant <= "001";
    konst_1257_wire_constant <= "0";
    konst_1260_wire_constant <= "010";
    konst_1263_wire_constant <= "0";
    konst_1267_wire_constant <= "011";
    konst_1270_wire_constant <= "0";
    konst_1273_wire_constant <= "100";
    konst_1276_wire_constant <= "0";
    konst_1293_wire_constant <= "001";
    konst_1297_wire_constant <= "0000000000000000";
    konst_1300_wire_constant <= "010";
    konst_1304_wire_constant <= "0000000000000000";
    konst_1308_wire_constant <= "011";
    konst_1312_wire_constant <= "0000000000000000";
    konst_1315_wire_constant <= "100";
    konst_1319_wire_constant <= "0000000000000000";
    konst_1326_wire_constant <= "000";
    konst_1329_wire_constant <= "0000000000000000";
    konst_1336_wire_constant <= "0000000000000001";
    konst_1340_wire_constant <= "0000000000000001";
    konst_1350_wire_constant <= "001";
    konst_1358_wire_constant <= "010";
    konst_1366_wire_constant <= "011";
    konst_1374_wire_constant <= "100";
    konst_1380_wire_constant <= "001";
    konst_1385_wire_constant <= "010";
    konst_1390_wire_constant <= "011";
    konst_1402_wire_constant <= "001";
    konst_1405_wire_constant <= "0";
    konst_1408_wire_constant <= "010";
    konst_1411_wire_constant <= "0";
    konst_1415_wire_constant <= "011";
    konst_1418_wire_constant <= "0";
    konst_1421_wire_constant <= "100";
    konst_1424_wire_constant <= "0";
    konst_1443_wire_constant <= "1";
    phi_stmt_1187: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1189_wire_constant & RPIPE_noblock_obuf_1_3_1191_wire;
      req <= phi_stmt_1187_req_0 & phi_stmt_1187_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1187",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1187_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1187,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1187
    phi_stmt_1192: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1194_wire_constant & RPIPE_noblock_obuf_2_3_1196_wire;
      req <= phi_stmt_1192_req_0 & phi_stmt_1192_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1192",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1192_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1192,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1192
    phi_stmt_1197: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1199_wire_constant & RPIPE_noblock_obuf_3_3_1201_wire;
      req <= phi_stmt_1197_req_0 & phi_stmt_1197_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1197",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1197_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1197,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1197
    phi_stmt_1202: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1204_wire_constant & RPIPE_noblock_obuf_4_3_1206_wire;
      req <= phi_stmt_1202_req_0 & phi_stmt_1202_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1202",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1202_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1202,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1202
    phi_stmt_1207: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1209_wire_constant & next_active_packet_1290_1210_buffered;
      req <= phi_stmt_1207_req_0 & phi_stmt_1207_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1207",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1207_ack_0,
          idata => idata,
          odata => active_packet_1207,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1207
    phi_stmt_1211: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_16_1213_wire_constant & next_down_counter_1345_1214_buffered;
      req <= phi_stmt_1211_req_0 & phi_stmt_1211_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1211",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1211_ack_0,
          idata => idata,
          odata => down_counter_1211,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1211
    phi_stmt_1215: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_1217_wire_constant & next_pkt_with_priority_1290_1218_buffered;
      req <= phi_stmt_1215_req_0 & phi_stmt_1215_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1215",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1215_ack_0,
          idata => idata,
          odata => pkt_with_priority_1215,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1215
    -- flow-through select operator MUX_1258_inst
    MUX_1258_wire <= p1_valid_1224 when (EQ_u3_u1_1255_wire(0) /=  '0') else konst_1257_wire_constant;
    -- flow-through select operator MUX_1264_inst
    MUX_1264_wire <= p2_valid_1229 when (EQ_u3_u1_1261_wire(0) /=  '0') else konst_1263_wire_constant;
    -- flow-through select operator MUX_1271_inst
    MUX_1271_wire <= p3_valid_1234 when (EQ_u3_u1_1268_wire(0) /=  '0') else konst_1270_wire_constant;
    -- flow-through select operator MUX_1277_inst
    MUX_1277_wire <= p4_valid_1239 when (EQ_u3_u1_1274_wire(0) /=  '0') else konst_1276_wire_constant;
    -- flow-through select operator MUX_1298_inst
    MUX_1298_wire <= slice_1296_wire when (EQ_u3_u1_1294_wire(0) /=  '0') else konst_1297_wire_constant;
    -- flow-through select operator MUX_1305_inst
    MUX_1305_wire <= slice_1303_wire when (EQ_u3_u1_1301_wire(0) /=  '0') else konst_1304_wire_constant;
    -- flow-through select operator MUX_1313_inst
    MUX_1313_wire <= slice_1311_wire when (EQ_u3_u1_1309_wire(0) /=  '0') else konst_1312_wire_constant;
    -- flow-through select operator MUX_1320_inst
    MUX_1320_wire <= slice_1318_wire when (EQ_u3_u1_1316_wire(0) /=  '0') else konst_1319_wire_constant;
    -- flow-through select operator MUX_1343_inst
    MUX_1343_wire <= SUB_u16_u16_1341_wire when (valid_active_pkt_word_read_1280(0) /=  '0') else down_counter_1211;
    -- flow-through select operator MUX_1344_inst
    next_down_counter_1345 <= SUB_u16_u16_1337_wire when (started_new_packet_1332(0) /=  '0') else MUX_1343_wire;
    -- flow-through select operator MUX_1396_inst
    MUX_1396_wire <= slice_1393_wire when (EQ_u3_u1_1391_wire(0) /=  '0') else slice_1395_wire;
    -- flow-through select operator MUX_1397_inst
    MUX_1397_wire <= slice_1388_wire when (EQ_u3_u1_1386_wire(0) /=  '0') else MUX_1396_wire;
    -- flow-through select operator MUX_1398_inst
    data_to_out_1399 <= slice_1383_wire when (EQ_u3_u1_1381_wire(0) /=  '0') else MUX_1397_wire;
    -- flow-through select operator MUX_1406_inst
    MUX_1406_wire <= p1_valid_1224 when (EQ_u3_u1_1403_wire(0) /=  '0') else konst_1405_wire_constant;
    -- flow-through select operator MUX_1412_inst
    MUX_1412_wire <= p2_valid_1229 when (EQ_u3_u1_1409_wire(0) /=  '0') else konst_1411_wire_constant;
    -- flow-through select operator MUX_1419_inst
    MUX_1419_wire <= p3_valid_1234 when (EQ_u3_u1_1416_wire(0) /=  '0') else konst_1418_wire_constant;
    -- flow-through select operator MUX_1425_inst
    MUX_1425_wire <= p4_valid_1239 when (EQ_u3_u1_1422_wire(0) /=  '0') else konst_1424_wire_constant;
    -- flow-through slice operator slice_1296_inst
    slice_1296_wire <= pkt_1_e_word_1187(23 downto 8);
    -- flow-through slice operator slice_1303_inst
    slice_1303_wire <= pkt_2_e_word_1192(23 downto 8);
    -- flow-through slice operator slice_1311_inst
    slice_1311_wire <= pkt_3_e_word_1197(23 downto 8);
    -- flow-through slice operator slice_1318_inst
    slice_1318_wire <= pkt_4_e_word_1202(23 downto 8);
    -- flow-through slice operator slice_1383_inst
    slice_1383_wire <= pkt_1_e_word_1187(31 downto 0);
    -- flow-through slice operator slice_1388_inst
    slice_1388_wire <= pkt_2_e_word_1192(31 downto 0);
    -- flow-through slice operator slice_1393_inst
    slice_1393_wire <= pkt_3_e_word_1197(31 downto 0);
    -- flow-through slice operator slice_1395_inst
    slice_1395_wire <= pkt_4_e_word_1202(31 downto 0);
    next_active_packet_1290_1210_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1290_1210_buf_req_0;
      next_active_packet_1290_1210_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1290_1210_buf_req_1;
      next_active_packet_1290_1210_buf_ack_1<= rack(0);
      next_active_packet_1290_1210_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1290_1210_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1290_1210_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1345_1214_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1345_1214_buf_req_0;
      next_down_counter_1345_1214_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1345_1214_buf_req_1;
      next_down_counter_1345_1214_buf_ack_1<= rack(0);
      next_down_counter_1345_1214_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1345_1214_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1345,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1345_1214_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_with_priority_1290_1218_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_with_priority_1290_1218_buf_req_0;
      next_pkt_with_priority_1290_1218_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_with_priority_1290_1218_buf_req_1;
      next_pkt_with_priority_1290_1218_buf_ack_1<= rack(0);
      next_pkt_with_priority_1290_1218_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_with_priority_1290_1218_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_with_priority_1290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_with_priority_1290_1218_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1185_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1443_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1185_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1185_branch_req_0,
          ack0 => do_while_stmt_1185_branch_ack_0,
          ack1 => do_while_stmt_1185_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1331_inst
    process(NEQ_u3_u1_1327_wire, EQ_u16_u1_1330_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u3_u1_1327_wire, EQ_u16_u1_1330_wire, tmp_var);
      started_new_packet_1332 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1223_inst
    process(pkt_1_e_word_1187) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1187, konst_1222_wire_constant, tmp_var);
      p1_valid_1224 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1228_inst
    process(pkt_2_e_word_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1192, konst_1227_wire_constant, tmp_var);
      p2_valid_1229 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1233_inst
    process(pkt_3_e_word_1197) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1197, konst_1232_wire_constant, tmp_var);
      p3_valid_1234 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1238_inst
    process(pkt_4_e_word_1202) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1202, konst_1237_wire_constant, tmp_var);
      p4_valid_1239 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1330_inst
    process(down_counter_1211) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1211, konst_1329_wire_constant, tmp_var);
      EQ_u16_u1_1330_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1255_inst
    process(active_packet_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1207, konst_1254_wire_constant, tmp_var);
      EQ_u3_u1_1255_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1261_inst
    process(active_packet_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1207, konst_1260_wire_constant, tmp_var);
      EQ_u3_u1_1261_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1268_inst
    process(active_packet_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1207, konst_1267_wire_constant, tmp_var);
      EQ_u3_u1_1268_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1274_inst
    process(active_packet_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1207, konst_1273_wire_constant, tmp_var);
      EQ_u3_u1_1274_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1294_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1293_wire_constant, tmp_var);
      EQ_u3_u1_1294_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1301_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1300_wire_constant, tmp_var);
      EQ_u3_u1_1301_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1309_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1308_wire_constant, tmp_var);
      EQ_u3_u1_1309_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1316_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1315_wire_constant, tmp_var);
      EQ_u3_u1_1316_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1351_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1350_wire_constant, tmp_var);
      EQ_u3_u1_1351_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1359_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1358_wire_constant, tmp_var);
      EQ_u3_u1_1359_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1367_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1366_wire_constant, tmp_var);
      EQ_u3_u1_1367_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1375_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1374_wire_constant, tmp_var);
      EQ_u3_u1_1375_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1381_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1380_wire_constant, tmp_var);
      EQ_u3_u1_1381_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1386_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1385_wire_constant, tmp_var);
      EQ_u3_u1_1386_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1391_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1390_wire_constant, tmp_var);
      EQ_u3_u1_1391_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1403_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1402_wire_constant, tmp_var);
      EQ_u3_u1_1403_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1409_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1408_wire_constant, tmp_var);
      EQ_u3_u1_1409_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1416_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1415_wire_constant, tmp_var);
      EQ_u3_u1_1416_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1422_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1290, konst_1421_wire_constant, tmp_var);
      EQ_u3_u1_1422_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_1327_inst
    process(next_active_packet_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_1290, konst_1326_wire_constant, tmp_var);
      NEQ_u3_u1_1327_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1348_inst
    process(p1_valid_1224) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1224, tmp_var);
      NOT_u1_u1_1348_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1356_inst
    process(p2_valid_1229) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1229, tmp_var);
      NOT_u1_u1_1356_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1364_inst
    process(p3_valid_1234) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1234, tmp_var);
      NOT_u1_u1_1364_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1372_inst
    process(p4_valid_1239) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1239, tmp_var);
      NOT_u1_u1_1372_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_1306_inst
    process(MUX_1298_wire, MUX_1305_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1298_wire, MUX_1305_wire, tmp_var);
      OR_u16_u16_1306_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1321_inst
    process(MUX_1313_wire, MUX_1320_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1313_wire, MUX_1320_wire, tmp_var);
      OR_u16_u16_1321_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1322_inst
    process(OR_u16_u16_1306_wire, OR_u16_u16_1321_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u16_u16_1306_wire, OR_u16_u16_1321_wire, tmp_var);
      valid_active_pkt_length_1323 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1265_inst
    process(MUX_1258_wire, MUX_1264_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1258_wire, MUX_1264_wire, tmp_var);
      OR_u1_u1_1265_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1278_inst
    process(MUX_1271_wire, MUX_1277_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1271_wire, MUX_1277_wire, tmp_var);
      OR_u1_u1_1278_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1279_inst
    process(OR_u1_u1_1265_wire, OR_u1_u1_1278_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1265_wire, OR_u1_u1_1278_wire, tmp_var);
      valid_active_pkt_word_read_1280 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1352_inst
    process(NOT_u1_u1_1348_wire, EQ_u3_u1_1351_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1348_wire, EQ_u3_u1_1351_wire, tmp_var);
      read_from_1_1353 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1360_inst
    process(NOT_u1_u1_1356_wire, EQ_u3_u1_1359_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1356_wire, EQ_u3_u1_1359_wire, tmp_var);
      read_from_2_1361 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1368_inst
    process(NOT_u1_u1_1364_wire, EQ_u3_u1_1367_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1364_wire, EQ_u3_u1_1367_wire, tmp_var);
      read_from_3_1369 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1376_inst
    process(NOT_u1_u1_1372_wire, EQ_u3_u1_1375_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1372_wire, EQ_u3_u1_1375_wire, tmp_var);
      read_from_4_1377 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1413_inst
    process(MUX_1406_wire, MUX_1412_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1406_wire, MUX_1412_wire, tmp_var);
      OR_u1_u1_1413_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1426_inst
    process(MUX_1419_wire, MUX_1425_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1419_wire, MUX_1425_wire, tmp_var);
      OR_u1_u1_1426_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1427_inst
    process(OR_u1_u1_1413_wire, OR_u1_u1_1426_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1413_wire, OR_u1_u1_1426_wire, tmp_var);
      send_flag_1428 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1337_inst
    process(valid_active_pkt_length_1323) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(valid_active_pkt_length_1323, konst_1336_wire_constant, tmp_var);
      SUB_u16_u16_1337_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1341_inst
    process(down_counter_1211) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_1211, konst_1340_wire_constant, tmp_var);
      SUB_u16_u16_1341_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_3_1191_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_3_1191_inst_req_0;
      RPIPE_noblock_obuf_1_3_1191_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_3_1191_inst_req_1;
      RPIPE_noblock_obuf_1_3_1191_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1353(0);
      RPIPE_noblock_obuf_1_3_1191_wire <= data_out(32 downto 0);
      noblock_obuf_1_3_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_3_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_3_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_3_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_3_pipe_read_req(0),
          oack => noblock_obuf_1_3_pipe_read_ack(0),
          odata => noblock_obuf_1_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_3_1196_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_3_1196_inst_req_0;
      RPIPE_noblock_obuf_2_3_1196_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_3_1196_inst_req_1;
      RPIPE_noblock_obuf_2_3_1196_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1361(0);
      RPIPE_noblock_obuf_2_3_1196_wire <= data_out(32 downto 0);
      noblock_obuf_2_3_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_3_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_3_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_3_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_3_pipe_read_req(0),
          oack => noblock_obuf_2_3_pipe_read_ack(0),
          odata => noblock_obuf_2_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_3_1201_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_3_1201_inst_req_0;
      RPIPE_noblock_obuf_3_3_1201_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_3_1201_inst_req_1;
      RPIPE_noblock_obuf_3_3_1201_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1369(0);
      RPIPE_noblock_obuf_3_3_1201_wire <= data_out(32 downto 0);
      noblock_obuf_3_3_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_3_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_3_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_3_pipe_read_req(0),
          oack => noblock_obuf_3_3_pipe_read_ack(0),
          odata => noblock_obuf_3_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_3_1206_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_3_1206_inst_req_0;
      RPIPE_noblock_obuf_4_3_1206_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_3_1206_inst_req_1;
      RPIPE_noblock_obuf_4_3_1206_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1377(0);
      RPIPE_noblock_obuf_4_3_1206_wire <= data_out(32 downto 0);
      noblock_obuf_4_3_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_3_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_3_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_3_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_3_pipe_read_req(0),
          oack => noblock_obuf_4_3_pipe_read_ack(0),
          odata => noblock_obuf_4_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_3_1430_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_3_1430_inst_req_0;
      WPIPE_out_data_3_1430_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_3_1430_inst_req_1;
      WPIPE_out_data_3_1430_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1428(0);
      data_in <= data_to_out_1399;
      out_data_3_write_0_gI: SplitGuardInterface generic map(name => "out_data_3_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_3_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_3", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_3_pipe_write_req(0),
          oack => out_data_3_pipe_write_ack(0),
          odata => out_data_3_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_3155: prioritySelect_Volatile port map(down_counter => down_counter_1211, active_packet => active_packet_1207, pkt_with_priority => pkt_with_priority_1215, p1_valid => p1_valid_1224, p2_valid => p2_valid_1229, p3_valid => p3_valid_1234, p4_valid => p4_valid_1239, next_active_packet => next_active_packet_1290, next_pkt_with_priority => next_pkt_with_priority_1290); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_3_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_4_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_4_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_4_Daemon;
architecture outputPort_4_Daemon_arch of outputPort_4_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_4_Daemon_CP_1900_start: Boolean;
  signal outputPort_4_Daemon_CP_1900_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(15 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_with_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_with_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal RPIPE_noblock_obuf_3_4_1464_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_3_4_1464_inst_req_0 : boolean;
  signal phi_stmt_1465_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_4_1454_inst_ack_1 : boolean;
  signal phi_stmt_1460_ack_0 : boolean;
  signal phi_stmt_1460_req_0 : boolean;
  signal phi_stmt_1465_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1454_inst_req_1 : boolean;
  signal phi_stmt_1455_req_1 : boolean;
  signal phi_stmt_1460_req_1 : boolean;
  signal phi_stmt_1455_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_4_1459_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_4_1459_inst_ack_0 : boolean;
  signal phi_stmt_1455_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1454_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_4_1464_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1454_inst_req_0 : boolean;
  signal phi_stmt_1465_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_4_1459_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_4_1464_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1459_inst_ack_1 : boolean;
  signal next_active_packet_1553_1473_buf_ack_0 : boolean;
  signal next_active_packet_1553_1473_buf_ack_1 : boolean;
  signal next_active_packet_1553_1473_buf_req_1 : boolean;
  signal phi_stmt_1470_ack_0 : boolean;
  signal phi_stmt_1470_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1469_inst_ack_1 : boolean;
  signal phi_stmt_1470_req_1 : boolean;
  signal next_active_packet_1553_1473_buf_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1469_inst_req_1 : boolean;
  signal phi_stmt_1474_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_4_1469_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1469_inst_req_0 : boolean;
  signal do_while_stmt_1448_branch_req_0 : boolean;
  signal phi_stmt_1450_req_1 : boolean;
  signal phi_stmt_1450_req_0 : boolean;
  signal phi_stmt_1450_ack_0 : boolean;
  signal phi_stmt_1474_req_0 : boolean;
  signal phi_stmt_1474_ack_0 : boolean;
  signal next_down_counter_1608_1477_buf_req_0 : boolean;
  signal next_down_counter_1608_1477_buf_ack_0 : boolean;
  signal next_down_counter_1608_1477_buf_req_1 : boolean;
  signal next_down_counter_1608_1477_buf_ack_1 : boolean;
  signal phi_stmt_1478_req_1 : boolean;
  signal phi_stmt_1478_req_0 : boolean;
  signal phi_stmt_1478_ack_0 : boolean;
  signal next_pkt_with_priority_1553_1481_buf_req_0 : boolean;
  signal next_pkt_with_priority_1553_1481_buf_ack_0 : boolean;
  signal next_pkt_with_priority_1553_1481_buf_req_1 : boolean;
  signal next_pkt_with_priority_1553_1481_buf_ack_1 : boolean;
  signal WPIPE_out_data_4_1693_inst_req_0 : boolean;
  signal WPIPE_out_data_4_1693_inst_ack_0 : boolean;
  signal WPIPE_out_data_4_1693_inst_req_1 : boolean;
  signal WPIPE_out_data_4_1693_inst_ack_1 : boolean;
  signal do_while_stmt_1448_branch_ack_0 : boolean;
  signal do_while_stmt_1448_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_4_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_4_Daemon_CP_1900_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_4_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_4_Daemon_CP_1900: Block -- control-path 
    signal outputPort_4_Daemon_CP_1900_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_4_Daemon_CP_1900_elements(0) <= outputPort_4_Daemon_CP_1900_start;
    outputPort_4_Daemon_CP_1900_symbol <= outputPort_4_Daemon_CP_1900_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1447/$entry
      -- CP-element group 0: 	 branch_block_stmt_1447/branch_block_stmt_1447__entry__
      -- CP-element group 0: 	 branch_block_stmt_1447/do_while_stmt_1448__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1447/$exit
      -- CP-element group 1: 	 branch_block_stmt_1447/branch_block_stmt_1447__exit__
      -- CP-element group 1: 	 branch_block_stmt_1447/do_while_stmt_1448__exit__
      -- 
    outputPort_4_Daemon_CP_1900_elements(1) <= outputPort_4_Daemon_CP_1900_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1447/do_while_stmt_1448/$entry
      -- CP-element group 2: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448__entry__
      -- 
    outputPort_4_Daemon_CP_1900_elements(2) <= outputPort_4_Daemon_CP_1900_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448__exit__
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1447/do_while_stmt_1448/loop_back
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	160 
    -- CP-element group 5: 	159 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1447/do_while_stmt_1448/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1447/do_while_stmt_1448/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1447/do_while_stmt_1448/loop_taken/$entry
      -- 
    outputPort_4_Daemon_CP_1900_elements(5) <= outputPort_4_Daemon_CP_1900_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1447/do_while_stmt_1448/loop_body_done
      -- 
    outputPort_4_Daemon_CP_1900_elements(6) <= outputPort_4_Daemon_CP_1900_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	42 
    -- CP-element group 7: 	63 
    -- CP-element group 7: 	84 
    -- CP-element group 7: 	105 
    -- CP-element group 7: 	124 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/back_edge_to_loop_body
      -- 
    outputPort_4_Daemon_CP_1900_elements(7) <= outputPort_4_Daemon_CP_1900_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	44 
    -- CP-element group 8: 	65 
    -- CP-element group 8: 	86 
    -- CP-element group 8: 	107 
    -- CP-element group 8: 	126 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/first_time_through_loop_body
      -- 
    outputPort_4_Daemon_CP_1900_elements(8) <= outputPort_4_Daemon_CP_1900_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	57 
    -- CP-element group 9: 	58 
    -- CP-element group 9: 	78 
    -- CP-element group 9: 	79 
    -- CP-element group 9: 	99 
    -- CP-element group 9: 	100 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	138 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/loop_body_start
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/condition_evaluated
      -- 
    condition_evaluated_1924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(10), ack => do_while_stmt_1448_branch_req_0); -- 
    outputPort_4_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(157) & outputPort_4_Daemon_CP_1900_elements(14);
      gj_outputPort_4_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11: 	99 
    -- CP-element group 11: 	118 
    -- CP-element group 11: 	137 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	38 
    -- CP-element group 11: 	59 
    -- CP-element group 11: 	80 
    -- CP-element group 11: 	101 
    -- CP-element group 11: 	120 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_sample_start__ps
      -- 
    outputPort_4_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(15) & outputPort_4_Daemon_CP_1900_elements(36) & outputPort_4_Daemon_CP_1900_elements(57) & outputPort_4_Daemon_CP_1900_elements(78) & outputPort_4_Daemon_CP_1900_elements(99) & outputPort_4_Daemon_CP_1900_elements(118) & outputPort_4_Daemon_CP_1900_elements(137) & outputPort_4_Daemon_CP_1900_elements(14);
      gj_outputPort_4_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	139 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	39 
    -- CP-element group 12: 	60 
    -- CP-element group 12: 	81 
    -- CP-element group 12: 	102 
    -- CP-element group 12: 	121 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	57 
    -- CP-element group 12: 	78 
    -- CP-element group 12: 	99 
    -- CP-element group 12: 	118 
    -- CP-element group 12: 	137 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_sample_completed_
      -- 
    outputPort_4_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(139) & outputPort_4_Daemon_CP_1900_elements(18) & outputPort_4_Daemon_CP_1900_elements(39) & outputPort_4_Daemon_CP_1900_elements(60) & outputPort_4_Daemon_CP_1900_elements(81) & outputPort_4_Daemon_CP_1900_elements(102) & outputPort_4_Daemon_CP_1900_elements(121);
      gj_outputPort_4_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	58 
    -- CP-element group 13: 	79 
    -- CP-element group 13: 	100 
    -- CP-element group 13: 	119 
    -- CP-element group 13: 	138 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	40 
    -- CP-element group 13: 	61 
    -- CP-element group 13: 	82 
    -- CP-element group 13: 	103 
    -- CP-element group 13: 	122 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_update_start__ps
      -- 
    outputPort_4_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(16) & outputPort_4_Daemon_CP_1900_elements(37) & outputPort_4_Daemon_CP_1900_elements(58) & outputPort_4_Daemon_CP_1900_elements(79) & outputPort_4_Daemon_CP_1900_elements(100) & outputPort_4_Daemon_CP_1900_elements(119) & outputPort_4_Daemon_CP_1900_elements(138);
      gj_outputPort_4_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	41 
    -- CP-element group 14: 	62 
    -- CP-element group 14: 	83 
    -- CP-element group 14: 	104 
    -- CP-element group 14: 	123 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_4_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(140) & outputPort_4_Daemon_CP_1900_elements(20) & outputPort_4_Daemon_CP_1900_elements(41) & outputPort_4_Daemon_CP_1900_elements(62) & outputPort_4_Daemon_CP_1900_elements(83) & outputPort_4_Daemon_CP_1900_elements(104) & outputPort_4_Daemon_CP_1900_elements(123);
      gj_outputPort_4_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(17) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(19) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(21) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_loopback_sample_req_ps
      -- 
    phi_stmt_1450_loopback_sample_req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1450_loopback_sample_req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(22), ack => phi_stmt_1450_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(23) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_entry_sample_req_ps
      -- 
    phi_stmt_1450_entry_sample_req_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1450_entry_sample_req_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(24), ack => phi_stmt_1450_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1450_phi_mux_ack_ps
      -- 
    phi_stmt_1450_phi_mux_ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1450_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1452_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1452_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1452_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1452_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1452_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1452_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1452_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(28) <= outputPort_4_Daemon_CP_1900_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1452_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(27), ack => outputPort_4_Daemon_CP_1900_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	35 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_Sample/$entry
      -- 
    rr_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(32), ack => RPIPE_noblock_obuf_1_4_1454_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(30) & outputPort_4_Daemon_CP_1900_elements(35);
      gj_outputPort_4_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: 	34 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_update_start_
      -- 
    cr_1971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(33), ack => RPIPE_noblock_obuf_1_4_1454_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(31) & outputPort_4_Daemon_CP_1900_elements(34);
      gj_outputPort_4_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	33 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_Sample/$exit
      -- 
    ra_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_4_1454_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	32 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_1_4_1454_update_completed_
      -- 
    ca_1972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_4_1454_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	11 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	155 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	11 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(38) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	12 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	13 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(40) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	154 
    -- CP-element group 41: 	14 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_update_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	7 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(42) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_loopback_sample_req_ps
      -- 
    phi_stmt_1455_loopback_sample_req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1455_loopback_sample_req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(43), ack => phi_stmt_1455_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	8 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(44) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_entry_sample_req
      -- CP-element group 45: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_entry_sample_req_ps
      -- 
    phi_stmt_1455_entry_sample_req_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1455_entry_sample_req_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(45), ack => phi_stmt_1455_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_phi_mux_ack_ps
      -- CP-element group 46: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1455_phi_mux_ack
      -- 
    phi_stmt_1455_phi_mux_ack_1989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1455_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1457_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1457_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1457_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1457_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1457_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1457_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1457_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(49) <= outputPort_4_Daemon_CP_1900_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1457_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(48), ack => outputPort_4_Daemon_CP_1900_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	56 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_Sample/rr
      -- 
    rr_2010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(53), ack => RPIPE_noblock_obuf_2_4_1459_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(51) & outputPort_4_Daemon_CP_1900_elements(56);
      gj_outputPort_4_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: 	55 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_Update/cr
      -- 
    cr_2015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(54), ack => RPIPE_noblock_obuf_2_4_1459_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(52) & outputPort_4_Daemon_CP_1900_elements(55);
      gj_outputPort_4_Daemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	54 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_Sample/ra
      -- 
    ra_2011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_4_1459_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	53 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_2_4_1459_Update/ca
      -- 
    ca_2016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_4_1459_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(56)); -- 
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	9 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	12 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	11 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	9 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	155 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	13 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	11 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(59) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	12 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	13 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(61) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	154 
    -- CP-element group 62: 	14 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_update_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	7 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(63) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_loopback_sample_req
      -- CP-element group 64: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_loopback_sample_req_ps
      -- 
    phi_stmt_1460_loopback_sample_req_2027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1460_loopback_sample_req_2027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(64), ack => phi_stmt_1460_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	8 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(65) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_entry_sample_req_ps
      -- CP-element group 66: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_entry_sample_req
      -- 
    phi_stmt_1460_entry_sample_req_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1460_entry_sample_req_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(66), ack => phi_stmt_1460_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_phi_mux_ack_ps
      -- CP-element group 67: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1460_phi_mux_ack
      -- 
    phi_stmt_1460_phi_mux_ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1460_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1462_sample_start__ps
      -- CP-element group 68: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1462_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1462_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1462_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1462_update_start__ps
      -- CP-element group 69: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1462_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1462_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(70) <= outputPort_4_Daemon_CP_1900_elements(71);
    -- CP-element group 71:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	70 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1462_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(69), ack => outputPort_4_Daemon_CP_1900_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	77 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_sample_start_
      -- 
    rr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(74), ack => RPIPE_noblock_obuf_3_4_1464_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(72) & outputPort_4_Daemon_CP_1900_elements(77);
      gj_outputPort_4_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	76 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_Update/cr
      -- 
    cr_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(75), ack => RPIPE_noblock_obuf_3_4_1464_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(73) & outputPort_4_Daemon_CP_1900_elements(76);
      gj_outputPort_4_Daemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	75 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_Sample/ra
      -- 
    ra_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_4_1464_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(76)); -- 
    -- CP-element group 77:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	74 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_3_4_1464_update_completed__ps
      -- 
    ca_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_4_1464_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	12 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	11 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	9 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	155 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	13 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	11 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(80) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 81:  join  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	12 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	13 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(82) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	154 
    -- CP-element group 83: 	14 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	7 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(84) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_loopback_sample_req
      -- CP-element group 85: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_loopback_sample_req_ps
      -- 
    phi_stmt_1465_loopback_sample_req_2071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1465_loopback_sample_req_2071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(85), ack => phi_stmt_1465_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	8 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(86) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 87:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_entry_sample_req
      -- CP-element group 87: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_entry_sample_req_ps
      -- 
    phi_stmt_1465_entry_sample_req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1465_entry_sample_req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(87), ack => phi_stmt_1465_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_phi_mux_ack_ps
      -- CP-element group 88: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1465_phi_mux_ack
      -- 
    phi_stmt_1465_phi_mux_ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1465_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1467_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1467_sample_start__ps
      -- CP-element group 89: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1467_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1467_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1467_update_start__ps
      -- CP-element group 90: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1467_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1467_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(91) <= outputPort_4_Daemon_CP_1900_elements(92);
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_33_1467_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(90), ack => outputPort_4_Daemon_CP_1900_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	98 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_Sample/$entry
      -- 
    rr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(95), ack => RPIPE_noblock_obuf_4_4_1469_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(93) & outputPort_4_Daemon_CP_1900_elements(98);
      gj_outputPort_4_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	97 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_update_start_
      -- CP-element group 96: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_Update/cr
      -- 
    cr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(96), ack => RPIPE_noblock_obuf_4_4_1469_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(94) & outputPort_4_Daemon_CP_1900_elements(97);
      gj_outputPort_4_Daemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	96 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_sample_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_Sample/$exit
      -- 
    ra_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_4_1469_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(97)); -- 
    -- CP-element group 98:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	95 
    -- CP-element group 98:  members (4) 
      -- CP-element group 98: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_update_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/RPIPE_noblock_obuf_4_4_1469_Update/ca
      -- 
    ca_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_4_1469_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(98)); -- 
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	9 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	12 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	11 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	9 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	155 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	13 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	11 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(101) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	12 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	13 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(103) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	154 
    -- CP-element group 104: 	14 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	7 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(105) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_loopback_sample_req_ps
      -- CP-element group 106: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_loopback_sample_req
      -- 
    phi_stmt_1470_loopback_sample_req_2115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1470_loopback_sample_req_2115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(106), ack => phi_stmt_1470_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(106) is bound as output of CP function.
    -- CP-element group 107:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	8 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(107) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 108:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_entry_sample_req_ps
      -- CP-element group 108: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_entry_sample_req
      -- 
    phi_stmt_1470_entry_sample_req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1470_entry_sample_req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(108), ack => phi_stmt_1470_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_phi_mux_ack_ps
      -- CP-element group 109: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1470_phi_mux_ack
      -- 
    phi_stmt_1470_phi_mux_ack_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1470_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(109)); -- 
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (4) 
      -- CP-element group 110: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_3_1472_sample_completed__ps
      -- CP-element group 110: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_3_1472_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_3_1472_sample_start__ps
      -- CP-element group 110: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_3_1472_sample_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_3_1472_update_start__ps
      -- CP-element group 111: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_3_1472_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_3_1472_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(112) <= outputPort_4_Daemon_CP_1900_elements(113);
    -- CP-element group 113:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	112 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_3_1472_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(113) is a control-delay.
    cp_element_113_delay: control_delay_element  generic map(name => " 113_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(111), ack => outputPort_4_Daemon_CP_1900_elements(113), clk => clk, reset =>reset);
    -- CP-element group 114:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_Sample/req
      -- 
    req_2142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(114), ack => next_active_packet_1553_1473_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_Update/req
      -- CP-element group 115: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_update_start_
      -- 
    req_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(115), ack => next_active_packet_1553_1473_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_Sample/ack
      -- CP-element group 116: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_sample_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_sample_completed_
      -- 
    ack_2143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1553_1473_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(116)); -- 
    -- CP-element group 117:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_Update/ack
      -- CP-element group 117: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_active_packet_1473_update_completed__ps
      -- 
    ack_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1553_1473_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	12 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	11 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	155 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	13 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	11 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(120) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	12 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	13 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(122) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	154 
    -- CP-element group 123: 	14 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_update_completed__ps
      -- CP-element group 123: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	7 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(124) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_loopback_sample_req_ps
      -- CP-element group 125: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_loopback_sample_req
      -- 
    phi_stmt_1474_loopback_sample_req_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1474_loopback_sample_req_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(125), ack => phi_stmt_1474_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	8 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(126) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_entry_sample_req
      -- CP-element group 127: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_entry_sample_req_ps
      -- 
    phi_stmt_1474_entry_sample_req_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1474_entry_sample_req_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(127), ack => phi_stmt_1474_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_phi_mux_ack
      -- CP-element group 128: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1474_phi_mux_ack_ps
      -- 
    phi_stmt_1474_phi_mux_ack_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1474_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (4) 
      -- CP-element group 129: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_16_1476_sample_start__ps
      -- CP-element group 129: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_16_1476_sample_completed__ps
      -- CP-element group 129: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_16_1476_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_16_1476_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_16_1476_update_start__ps
      -- CP-element group 130: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_16_1476_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_16_1476_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(131) <= outputPort_4_Daemon_CP_1900_elements(132);
    -- CP-element group 132:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	131 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_ZERO_16_1476_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(132) is a control-delay.
    cp_element_132_delay: control_delay_element  generic map(name => " 132_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(130), ack => outputPort_4_Daemon_CP_1900_elements(132), clk => clk, reset =>reset);
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_Sample/req
      -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(133), ack => next_down_counter_1608_1477_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_update_start_
      -- CP-element group 134: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_Update/req
      -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(134), ack => next_down_counter_1608_1477_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_sample_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_Sample/ack
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1608_1477_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(135)); -- 
    -- CP-element group 136:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_update_completed__ps
      -- CP-element group 136: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_down_counter_1477_Update/ack
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1608_1477_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(136)); -- 
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	12 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	11 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	155 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	13 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	12 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(141) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_loopback_sample_req_ps
      -- 
    phi_stmt_1478_loopback_sample_req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1478_loopback_sample_req_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(142), ack => phi_stmt_1478_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(143) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_entry_sample_req_ps
      -- 
    phi_stmt_1478_entry_sample_req_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1478_entry_sample_req_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(144), ack => phi_stmt_1478_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/phi_stmt_1478_phi_mux_ack_ps
      -- 
    phi_stmt_1478_phi_mux_ack_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1478_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/konst_1480_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/konst_1480_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/konst_1480_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/konst_1480_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/konst_1480_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/konst_1480_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/konst_1480_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(148) <= outputPort_4_Daemon_CP_1900_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/konst_1480_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(147), ack => outputPort_4_Daemon_CP_1900_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_Sample/req
      -- 
    req_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(150), ack => next_pkt_with_priority_1553_1481_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_Update/req
      -- 
    req_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(151), ack => next_pkt_with_priority_1553_1481_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_Sample/ack
      -- 
    ack_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_with_priority_1553_1481_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/R_next_pkt_with_priority_1481_Update/ack
      -- 
    ack_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_with_priority_1553_1481_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	41 
    -- CP-element group 154: 	62 
    -- CP-element group 154: 	83 
    -- CP-element group 154: 	104 
    -- CP-element group 154: 	123 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_Sample/req
      -- 
    req_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(154), ack => WPIPE_out_data_4_1693_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(140) & outputPort_4_Daemon_CP_1900_elements(20) & outputPort_4_Daemon_CP_1900_elements(41) & outputPort_4_Daemon_CP_1900_elements(62) & outputPort_4_Daemon_CP_1900_elements(83) & outputPort_4_Daemon_CP_1900_elements(104) & outputPort_4_Daemon_CP_1900_elements(123) & outputPort_4_Daemon_CP_1900_elements(156);
      gj_outputPort_4_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	37 
    -- CP-element group 155: 	58 
    -- CP-element group 155: 	79 
    -- CP-element group 155: 	100 
    -- CP-element group 155: 	119 
    -- CP-element group 155: 	138 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_Update/req
      -- 
    ack_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4_1693_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(155)); -- 
    req_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(155), ack => WPIPE_out_data_4_1693_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/WPIPE_out_data_4_1693_Update/ack
      -- 
    ack_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4_1693_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(9), ack => outputPort_4_Daemon_CP_1900_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1447/do_while_stmt_1448/do_while_stmt_1448_loop_body/$exit
      -- 
    outputPort_4_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(156) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_1447/do_while_stmt_1448/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_1447/do_while_stmt_1448/loop_exit/ack
      -- 
    ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1448_branch_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1447/do_while_stmt_1448/loop_taken/$exit
      -- CP-element group 160: 	 branch_block_stmt_1447/do_while_stmt_1448/loop_taken/ack
      -- 
    ack_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1448_branch_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1447/do_while_stmt_1448/$exit
      -- 
    outputPort_4_Daemon_CP_1900_elements(161) <= outputPort_4_Daemon_CP_1900_elements(3);
    outputPort_4_Daemon_do_while_stmt_1448_terminator_2261: loop_terminator -- 
      generic map (name => " outputPort_4_Daemon_do_while_stmt_1448_terminator_2261", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_4_Daemon_CP_1900_elements(6),loop_continue => outputPort_4_Daemon_CP_1900_elements(160),loop_terminate => outputPort_4_Daemon_CP_1900_elements(159),loop_back => outputPort_4_Daemon_CP_1900_elements(4),loop_exit => outputPort_4_Daemon_CP_1900_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1450_phi_seq_1973_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(23);
      outputPort_4_Daemon_CP_1900_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(26);
      outputPort_4_Daemon_CP_1900_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(28);
      outputPort_4_Daemon_CP_1900_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(21);
      outputPort_4_Daemon_CP_1900_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(34);
      outputPort_4_Daemon_CP_1900_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(35);
      outputPort_4_Daemon_CP_1900_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1450_phi_seq_1973 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1450_phi_seq_1973") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(17), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(18), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(19), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(20), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1455_phi_seq_2017_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(44);
      outputPort_4_Daemon_CP_1900_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(47);
      outputPort_4_Daemon_CP_1900_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(49);
      outputPort_4_Daemon_CP_1900_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(42);
      outputPort_4_Daemon_CP_1900_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(55);
      outputPort_4_Daemon_CP_1900_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(56);
      outputPort_4_Daemon_CP_1900_elements(43) <= phi_mux_reqs(1);
      phi_stmt_1455_phi_seq_2017 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1455_phi_seq_2017") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(38), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(39), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(40), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(41), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1460_phi_seq_2061_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(65);
      outputPort_4_Daemon_CP_1900_elements(68)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(68);
      outputPort_4_Daemon_CP_1900_elements(69)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(70);
      outputPort_4_Daemon_CP_1900_elements(66) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(63);
      outputPort_4_Daemon_CP_1900_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(76);
      outputPort_4_Daemon_CP_1900_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(77);
      outputPort_4_Daemon_CP_1900_elements(64) <= phi_mux_reqs(1);
      phi_stmt_1460_phi_seq_2061 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1460_phi_seq_2061") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(59), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(60), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(61), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(62), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(67), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1465_phi_seq_2105_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(86);
      outputPort_4_Daemon_CP_1900_elements(89)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(89);
      outputPort_4_Daemon_CP_1900_elements(90)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(91);
      outputPort_4_Daemon_CP_1900_elements(87) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(84);
      outputPort_4_Daemon_CP_1900_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(97);
      outputPort_4_Daemon_CP_1900_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(98);
      outputPort_4_Daemon_CP_1900_elements(85) <= phi_mux_reqs(1);
      phi_stmt_1465_phi_seq_2105 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1465_phi_seq_2105") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(80), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(81), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(82), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(83), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(88), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1470_phi_seq_2149_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(107);
      outputPort_4_Daemon_CP_1900_elements(110)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(110);
      outputPort_4_Daemon_CP_1900_elements(111)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(112);
      outputPort_4_Daemon_CP_1900_elements(108) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(105);
      outputPort_4_Daemon_CP_1900_elements(114)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(116);
      outputPort_4_Daemon_CP_1900_elements(115)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(117);
      outputPort_4_Daemon_CP_1900_elements(106) <= phi_mux_reqs(1);
      phi_stmt_1470_phi_seq_2149 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1470_phi_seq_2149") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(101), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(102), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(103), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(104), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(109), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1474_phi_seq_2193_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(126);
      outputPort_4_Daemon_CP_1900_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(129);
      outputPort_4_Daemon_CP_1900_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(131);
      outputPort_4_Daemon_CP_1900_elements(127) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(124);
      outputPort_4_Daemon_CP_1900_elements(133)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(135);
      outputPort_4_Daemon_CP_1900_elements(134)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(136);
      outputPort_4_Daemon_CP_1900_elements(125) <= phi_mux_reqs(1);
      phi_stmt_1474_phi_seq_2193 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1474_phi_seq_2193") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(120), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(121), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(122), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(123), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1478_phi_seq_2237_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(143);
      outputPort_4_Daemon_CP_1900_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(146);
      outputPort_4_Daemon_CP_1900_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(148);
      outputPort_4_Daemon_CP_1900_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(141);
      outputPort_4_Daemon_CP_1900_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(152);
      outputPort_4_Daemon_CP_1900_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(153);
      outputPort_4_Daemon_CP_1900_elements(142) <= phi_mux_reqs(1);
      phi_stmt_1478_phi_seq_2237 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1478_phi_seq_2237") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(11), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(139), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(13), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(140), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1925_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_4_Daemon_CP_1900_elements(7);
        preds(1)  <= outputPort_4_Daemon_CP_1900_elements(8);
        entry_tmerge_1925 : transition_merge -- 
          generic map(name => " entry_tmerge_1925")
          port map (preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u16_u1_1593_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1518_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1524_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1531_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1537_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1557_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1564_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1572_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1579_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1614_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1622_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1630_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1638_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1644_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1649_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1654_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1666_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1672_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1679_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1685_wire : std_logic_vector(0 downto 0);
    signal MUX_1521_wire : std_logic_vector(0 downto 0);
    signal MUX_1527_wire : std_logic_vector(0 downto 0);
    signal MUX_1534_wire : std_logic_vector(0 downto 0);
    signal MUX_1540_wire : std_logic_vector(0 downto 0);
    signal MUX_1561_wire : std_logic_vector(15 downto 0);
    signal MUX_1568_wire : std_logic_vector(15 downto 0);
    signal MUX_1576_wire : std_logic_vector(15 downto 0);
    signal MUX_1583_wire : std_logic_vector(15 downto 0);
    signal MUX_1606_wire : std_logic_vector(15 downto 0);
    signal MUX_1659_wire : std_logic_vector(31 downto 0);
    signal MUX_1660_wire : std_logic_vector(31 downto 0);
    signal MUX_1669_wire : std_logic_vector(0 downto 0);
    signal MUX_1675_wire : std_logic_vector(0 downto 0);
    signal MUX_1682_wire : std_logic_vector(0 downto 0);
    signal MUX_1688_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_1590_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1611_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1619_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1627_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1635_wire : std_logic_vector(0 downto 0);
    signal OR_u16_u16_1569_wire : std_logic_vector(15 downto 0);
    signal OR_u16_u16_1584_wire : std_logic_vector(15 downto 0);
    signal OR_u1_u1_1528_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1541_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1676_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1689_wire : std_logic_vector(0 downto 0);
    signal RPIPE_noblock_obuf_1_4_1454_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_4_1459_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_4_1464_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_4_1469_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_16_1476_wire_constant : std_logic_vector(15 downto 0);
    signal R_ZERO_33_1452_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1457_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1462_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1467_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1472_wire_constant : std_logic_vector(2 downto 0);
    signal SUB_u16_u16_1600_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_1604_wire : std_logic_vector(15 downto 0);
    signal active_packet_1470 : std_logic_vector(2 downto 0);
    signal data_to_out_1662 : std_logic_vector(31 downto 0);
    signal down_counter_1474 : std_logic_vector(15 downto 0);
    signal konst_1480_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1485_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1490_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1495_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1500_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1517_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1520_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1523_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1526_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1530_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1533_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1536_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1539_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1556_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1560_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1563_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1567_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1571_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1575_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1578_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1582_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1589_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1592_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1599_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1603_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1613_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1621_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1629_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1637_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1643_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1648_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1653_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1665_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1668_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1671_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1674_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1678_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1681_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1684_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1687_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1706_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1553 : std_logic_vector(2 downto 0);
    signal next_active_packet_1553_1473_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_1608 : std_logic_vector(15 downto 0);
    signal next_down_counter_1608_1477_buffered : std_logic_vector(15 downto 0);
    signal next_pkt_with_priority_1553 : std_logic_vector(2 downto 0);
    signal next_pkt_with_priority_1553_1481_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_1487 : std_logic_vector(0 downto 0);
    signal p2_valid_1492 : std_logic_vector(0 downto 0);
    signal p3_valid_1497 : std_logic_vector(0 downto 0);
    signal p4_valid_1502 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1450 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1455 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1460 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1465 : std_logic_vector(32 downto 0);
    signal pkt_with_priority_1478 : std_logic_vector(2 downto 0);
    signal read_from_1_1616 : std_logic_vector(0 downto 0);
    signal read_from_2_1624 : std_logic_vector(0 downto 0);
    signal read_from_3_1632 : std_logic_vector(0 downto 0);
    signal read_from_4_1640 : std_logic_vector(0 downto 0);
    signal send_flag_1691 : std_logic_vector(0 downto 0);
    signal slice_1559_wire : std_logic_vector(15 downto 0);
    signal slice_1566_wire : std_logic_vector(15 downto 0);
    signal slice_1574_wire : std_logic_vector(15 downto 0);
    signal slice_1581_wire : std_logic_vector(15 downto 0);
    signal slice_1646_wire : std_logic_vector(31 downto 0);
    signal slice_1651_wire : std_logic_vector(31 downto 0);
    signal slice_1656_wire : std_logic_vector(31 downto 0);
    signal slice_1658_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1595 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_length_1586 : std_logic_vector(15 downto 0);
    signal valid_active_pkt_word_read_1543 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_16_1476_wire_constant <= "0000000000000000";
    R_ZERO_33_1452_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1457_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1462_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1467_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1472_wire_constant <= "000";
    konst_1480_wire_constant <= "001";
    konst_1485_wire_constant <= "000000000000000000000000000100000";
    konst_1490_wire_constant <= "000000000000000000000000000100000";
    konst_1495_wire_constant <= "000000000000000000000000000100000";
    konst_1500_wire_constant <= "000000000000000000000000000100000";
    konst_1517_wire_constant <= "001";
    konst_1520_wire_constant <= "0";
    konst_1523_wire_constant <= "010";
    konst_1526_wire_constant <= "0";
    konst_1530_wire_constant <= "011";
    konst_1533_wire_constant <= "0";
    konst_1536_wire_constant <= "100";
    konst_1539_wire_constant <= "0";
    konst_1556_wire_constant <= "001";
    konst_1560_wire_constant <= "0000000000000000";
    konst_1563_wire_constant <= "010";
    konst_1567_wire_constant <= "0000000000000000";
    konst_1571_wire_constant <= "011";
    konst_1575_wire_constant <= "0000000000000000";
    konst_1578_wire_constant <= "100";
    konst_1582_wire_constant <= "0000000000000000";
    konst_1589_wire_constant <= "000";
    konst_1592_wire_constant <= "0000000000000000";
    konst_1599_wire_constant <= "0000000000000001";
    konst_1603_wire_constant <= "0000000000000001";
    konst_1613_wire_constant <= "001";
    konst_1621_wire_constant <= "010";
    konst_1629_wire_constant <= "011";
    konst_1637_wire_constant <= "100";
    konst_1643_wire_constant <= "001";
    konst_1648_wire_constant <= "010";
    konst_1653_wire_constant <= "011";
    konst_1665_wire_constant <= "001";
    konst_1668_wire_constant <= "0";
    konst_1671_wire_constant <= "010";
    konst_1674_wire_constant <= "0";
    konst_1678_wire_constant <= "011";
    konst_1681_wire_constant <= "0";
    konst_1684_wire_constant <= "100";
    konst_1687_wire_constant <= "0";
    konst_1706_wire_constant <= "1";
    phi_stmt_1450: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1452_wire_constant & RPIPE_noblock_obuf_1_4_1454_wire;
      req <= phi_stmt_1450_req_0 & phi_stmt_1450_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1450",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1450_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1450,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1450
    phi_stmt_1455: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1457_wire_constant & RPIPE_noblock_obuf_2_4_1459_wire;
      req <= phi_stmt_1455_req_0 & phi_stmt_1455_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1455",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1455_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1455,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1455
    phi_stmt_1460: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1462_wire_constant & RPIPE_noblock_obuf_3_4_1464_wire;
      req <= phi_stmt_1460_req_0 & phi_stmt_1460_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1460",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1460_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1460,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1460
    phi_stmt_1465: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1467_wire_constant & RPIPE_noblock_obuf_4_4_1469_wire;
      req <= phi_stmt_1465_req_0 & phi_stmt_1465_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1465",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1465_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1465,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1465
    phi_stmt_1470: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1472_wire_constant & next_active_packet_1553_1473_buffered;
      req <= phi_stmt_1470_req_0 & phi_stmt_1470_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1470",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1470_ack_0,
          idata => idata,
          odata => active_packet_1470,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1470
    phi_stmt_1474: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_16_1476_wire_constant & next_down_counter_1608_1477_buffered;
      req <= phi_stmt_1474_req_0 & phi_stmt_1474_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1474",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1474_ack_0,
          idata => idata,
          odata => down_counter_1474,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1474
    phi_stmt_1478: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_1480_wire_constant & next_pkt_with_priority_1553_1481_buffered;
      req <= phi_stmt_1478_req_0 & phi_stmt_1478_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1478",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1478_ack_0,
          idata => idata,
          odata => pkt_with_priority_1478,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1478
    -- flow-through select operator MUX_1521_inst
    MUX_1521_wire <= p1_valid_1487 when (EQ_u3_u1_1518_wire(0) /=  '0') else konst_1520_wire_constant;
    -- flow-through select operator MUX_1527_inst
    MUX_1527_wire <= p2_valid_1492 when (EQ_u3_u1_1524_wire(0) /=  '0') else konst_1526_wire_constant;
    -- flow-through select operator MUX_1534_inst
    MUX_1534_wire <= p3_valid_1497 when (EQ_u3_u1_1531_wire(0) /=  '0') else konst_1533_wire_constant;
    -- flow-through select operator MUX_1540_inst
    MUX_1540_wire <= p4_valid_1502 when (EQ_u3_u1_1537_wire(0) /=  '0') else konst_1539_wire_constant;
    -- flow-through select operator MUX_1561_inst
    MUX_1561_wire <= slice_1559_wire when (EQ_u3_u1_1557_wire(0) /=  '0') else konst_1560_wire_constant;
    -- flow-through select operator MUX_1568_inst
    MUX_1568_wire <= slice_1566_wire when (EQ_u3_u1_1564_wire(0) /=  '0') else konst_1567_wire_constant;
    -- flow-through select operator MUX_1576_inst
    MUX_1576_wire <= slice_1574_wire when (EQ_u3_u1_1572_wire(0) /=  '0') else konst_1575_wire_constant;
    -- flow-through select operator MUX_1583_inst
    MUX_1583_wire <= slice_1581_wire when (EQ_u3_u1_1579_wire(0) /=  '0') else konst_1582_wire_constant;
    -- flow-through select operator MUX_1606_inst
    MUX_1606_wire <= SUB_u16_u16_1604_wire when (valid_active_pkt_word_read_1543(0) /=  '0') else down_counter_1474;
    -- flow-through select operator MUX_1607_inst
    next_down_counter_1608 <= SUB_u16_u16_1600_wire when (started_new_packet_1595(0) /=  '0') else MUX_1606_wire;
    -- flow-through select operator MUX_1659_inst
    MUX_1659_wire <= slice_1656_wire when (EQ_u3_u1_1654_wire(0) /=  '0') else slice_1658_wire;
    -- flow-through select operator MUX_1660_inst
    MUX_1660_wire <= slice_1651_wire when (EQ_u3_u1_1649_wire(0) /=  '0') else MUX_1659_wire;
    -- flow-through select operator MUX_1661_inst
    data_to_out_1662 <= slice_1646_wire when (EQ_u3_u1_1644_wire(0) /=  '0') else MUX_1660_wire;
    -- flow-through select operator MUX_1669_inst
    MUX_1669_wire <= p1_valid_1487 when (EQ_u3_u1_1666_wire(0) /=  '0') else konst_1668_wire_constant;
    -- flow-through select operator MUX_1675_inst
    MUX_1675_wire <= p2_valid_1492 when (EQ_u3_u1_1672_wire(0) /=  '0') else konst_1674_wire_constant;
    -- flow-through select operator MUX_1682_inst
    MUX_1682_wire <= p3_valid_1497 when (EQ_u3_u1_1679_wire(0) /=  '0') else konst_1681_wire_constant;
    -- flow-through select operator MUX_1688_inst
    MUX_1688_wire <= p4_valid_1502 when (EQ_u3_u1_1685_wire(0) /=  '0') else konst_1687_wire_constant;
    -- flow-through slice operator slice_1559_inst
    slice_1559_wire <= pkt_1_e_word_1450(23 downto 8);
    -- flow-through slice operator slice_1566_inst
    slice_1566_wire <= pkt_2_e_word_1455(23 downto 8);
    -- flow-through slice operator slice_1574_inst
    slice_1574_wire <= pkt_3_e_word_1460(23 downto 8);
    -- flow-through slice operator slice_1581_inst
    slice_1581_wire <= pkt_4_e_word_1465(23 downto 8);
    -- flow-through slice operator slice_1646_inst
    slice_1646_wire <= pkt_1_e_word_1450(31 downto 0);
    -- flow-through slice operator slice_1651_inst
    slice_1651_wire <= pkt_2_e_word_1455(31 downto 0);
    -- flow-through slice operator slice_1656_inst
    slice_1656_wire <= pkt_3_e_word_1460(31 downto 0);
    -- flow-through slice operator slice_1658_inst
    slice_1658_wire <= pkt_4_e_word_1465(31 downto 0);
    next_active_packet_1553_1473_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1553_1473_buf_req_0;
      next_active_packet_1553_1473_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1553_1473_buf_req_1;
      next_active_packet_1553_1473_buf_ack_1<= rack(0);
      next_active_packet_1553_1473_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1553_1473_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1553_1473_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1608_1477_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1608_1477_buf_req_0;
      next_down_counter_1608_1477_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1608_1477_buf_req_1;
      next_down_counter_1608_1477_buf_ack_1<= rack(0);
      next_down_counter_1608_1477_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1608_1477_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1608_1477_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_with_priority_1553_1481_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_with_priority_1553_1481_buf_req_0;
      next_pkt_with_priority_1553_1481_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_with_priority_1553_1481_buf_req_1;
      next_pkt_with_priority_1553_1481_buf_ack_1<= rack(0);
      next_pkt_with_priority_1553_1481_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_with_priority_1553_1481_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_with_priority_1553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_with_priority_1553_1481_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1448_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1706_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1448_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1448_branch_req_0,
          ack0 => do_while_stmt_1448_branch_ack_0,
          ack1 => do_while_stmt_1448_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1594_inst
    process(NEQ_u3_u1_1590_wire, EQ_u16_u1_1593_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u3_u1_1590_wire, EQ_u16_u1_1593_wire, tmp_var);
      started_new_packet_1595 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1486_inst
    process(pkt_1_e_word_1450) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1450, konst_1485_wire_constant, tmp_var);
      p1_valid_1487 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1491_inst
    process(pkt_2_e_word_1455) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1455, konst_1490_wire_constant, tmp_var);
      p2_valid_1492 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1496_inst
    process(pkt_3_e_word_1460) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1460, konst_1495_wire_constant, tmp_var);
      p3_valid_1497 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1501_inst
    process(pkt_4_e_word_1465) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1465, konst_1500_wire_constant, tmp_var);
      p4_valid_1502 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1593_inst
    process(down_counter_1474) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1474, konst_1592_wire_constant, tmp_var);
      EQ_u16_u1_1593_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1518_inst
    process(active_packet_1470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1470, konst_1517_wire_constant, tmp_var);
      EQ_u3_u1_1518_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1524_inst
    process(active_packet_1470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1470, konst_1523_wire_constant, tmp_var);
      EQ_u3_u1_1524_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1531_inst
    process(active_packet_1470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1470, konst_1530_wire_constant, tmp_var);
      EQ_u3_u1_1531_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1537_inst
    process(active_packet_1470) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1470, konst_1536_wire_constant, tmp_var);
      EQ_u3_u1_1537_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1557_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1556_wire_constant, tmp_var);
      EQ_u3_u1_1557_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1564_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1563_wire_constant, tmp_var);
      EQ_u3_u1_1564_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1572_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1571_wire_constant, tmp_var);
      EQ_u3_u1_1572_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1579_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1578_wire_constant, tmp_var);
      EQ_u3_u1_1579_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1614_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1613_wire_constant, tmp_var);
      EQ_u3_u1_1614_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1622_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1621_wire_constant, tmp_var);
      EQ_u3_u1_1622_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1630_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1629_wire_constant, tmp_var);
      EQ_u3_u1_1630_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1638_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1637_wire_constant, tmp_var);
      EQ_u3_u1_1638_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1644_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1643_wire_constant, tmp_var);
      EQ_u3_u1_1644_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1649_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1648_wire_constant, tmp_var);
      EQ_u3_u1_1649_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1654_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1653_wire_constant, tmp_var);
      EQ_u3_u1_1654_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1666_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1665_wire_constant, tmp_var);
      EQ_u3_u1_1666_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1672_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1671_wire_constant, tmp_var);
      EQ_u3_u1_1672_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1679_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1678_wire_constant, tmp_var);
      EQ_u3_u1_1679_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1685_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1553, konst_1684_wire_constant, tmp_var);
      EQ_u3_u1_1685_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_1590_inst
    process(next_active_packet_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_1553, konst_1589_wire_constant, tmp_var);
      NEQ_u3_u1_1590_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1611_inst
    process(p1_valid_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1487, tmp_var);
      NOT_u1_u1_1611_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1619_inst
    process(p2_valid_1492) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1492, tmp_var);
      NOT_u1_u1_1619_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1627_inst
    process(p3_valid_1497) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1497, tmp_var);
      NOT_u1_u1_1627_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1635_inst
    process(p4_valid_1502) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1502, tmp_var);
      NOT_u1_u1_1635_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_1569_inst
    process(MUX_1561_wire, MUX_1568_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1561_wire, MUX_1568_wire, tmp_var);
      OR_u16_u16_1569_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1584_inst
    process(MUX_1576_wire, MUX_1583_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1576_wire, MUX_1583_wire, tmp_var);
      OR_u16_u16_1584_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1585_inst
    process(OR_u16_u16_1569_wire, OR_u16_u16_1584_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u16_u16_1569_wire, OR_u16_u16_1584_wire, tmp_var);
      valid_active_pkt_length_1586 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1528_inst
    process(MUX_1521_wire, MUX_1527_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1521_wire, MUX_1527_wire, tmp_var);
      OR_u1_u1_1528_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1541_inst
    process(MUX_1534_wire, MUX_1540_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1534_wire, MUX_1540_wire, tmp_var);
      OR_u1_u1_1541_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1542_inst
    process(OR_u1_u1_1528_wire, OR_u1_u1_1541_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1528_wire, OR_u1_u1_1541_wire, tmp_var);
      valid_active_pkt_word_read_1543 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1615_inst
    process(NOT_u1_u1_1611_wire, EQ_u3_u1_1614_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1611_wire, EQ_u3_u1_1614_wire, tmp_var);
      read_from_1_1616 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1623_inst
    process(NOT_u1_u1_1619_wire, EQ_u3_u1_1622_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1619_wire, EQ_u3_u1_1622_wire, tmp_var);
      read_from_2_1624 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1631_inst
    process(NOT_u1_u1_1627_wire, EQ_u3_u1_1630_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1627_wire, EQ_u3_u1_1630_wire, tmp_var);
      read_from_3_1632 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1639_inst
    process(NOT_u1_u1_1635_wire, EQ_u3_u1_1638_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1635_wire, EQ_u3_u1_1638_wire, tmp_var);
      read_from_4_1640 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1676_inst
    process(MUX_1669_wire, MUX_1675_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1669_wire, MUX_1675_wire, tmp_var);
      OR_u1_u1_1676_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1689_inst
    process(MUX_1682_wire, MUX_1688_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1682_wire, MUX_1688_wire, tmp_var);
      OR_u1_u1_1689_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1690_inst
    process(OR_u1_u1_1676_wire, OR_u1_u1_1689_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1676_wire, OR_u1_u1_1689_wire, tmp_var);
      send_flag_1691 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1600_inst
    process(valid_active_pkt_length_1586) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(valid_active_pkt_length_1586, konst_1599_wire_constant, tmp_var);
      SUB_u16_u16_1600_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1604_inst
    process(down_counter_1474) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_1474, konst_1603_wire_constant, tmp_var);
      SUB_u16_u16_1604_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_4_1454_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_4_1454_inst_req_0;
      RPIPE_noblock_obuf_1_4_1454_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_4_1454_inst_req_1;
      RPIPE_noblock_obuf_1_4_1454_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1616(0);
      RPIPE_noblock_obuf_1_4_1454_wire <= data_out(32 downto 0);
      noblock_obuf_1_4_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_4_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_4_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_4_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_4_pipe_read_req(0),
          oack => noblock_obuf_1_4_pipe_read_ack(0),
          odata => noblock_obuf_1_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_4_1459_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_4_1459_inst_req_0;
      RPIPE_noblock_obuf_2_4_1459_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_4_1459_inst_req_1;
      RPIPE_noblock_obuf_2_4_1459_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1624(0);
      RPIPE_noblock_obuf_2_4_1459_wire <= data_out(32 downto 0);
      noblock_obuf_2_4_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_4_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_4_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_4_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_4_pipe_read_req(0),
          oack => noblock_obuf_2_4_pipe_read_ack(0),
          odata => noblock_obuf_2_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_4_1464_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_4_1464_inst_req_0;
      RPIPE_noblock_obuf_3_4_1464_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_4_1464_inst_req_1;
      RPIPE_noblock_obuf_3_4_1464_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1632(0);
      RPIPE_noblock_obuf_3_4_1464_wire <= data_out(32 downto 0);
      noblock_obuf_3_4_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_4_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_4_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_4_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_4_pipe_read_req(0),
          oack => noblock_obuf_3_4_pipe_read_ack(0),
          odata => noblock_obuf_3_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_4_1469_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_4_1469_inst_req_0;
      RPIPE_noblock_obuf_4_4_1469_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_4_1469_inst_req_1;
      RPIPE_noblock_obuf_4_4_1469_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1640(0);
      RPIPE_noblock_obuf_4_4_1469_wire <= data_out(32 downto 0);
      noblock_obuf_4_4_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_4_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_4_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_4_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_4_pipe_read_req(0),
          oack => noblock_obuf_4_4_pipe_read_ack(0),
          odata => noblock_obuf_4_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_4_1693_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_4_1693_inst_req_0;
      WPIPE_out_data_4_1693_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_4_1693_inst_req_1;
      WPIPE_out_data_4_1693_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1691(0);
      data_in <= data_to_out_1662;
      out_data_4_write_0_gI: SplitGuardInterface generic map(name => "out_data_4_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_4_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_4", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_4_pipe_write_req(0),
          oack => out_data_4_pipe_write_ack(0),
          odata => out_data_4_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_3786: prioritySelect_Volatile port map(down_counter => down_counter_1474, active_packet => active_packet_1470, pkt_with_priority => pkt_with_priority_1478, p1_valid => p1_valid_1487, p2_valid => p2_valid_1492, p3_valid => p3_valid_1497, p4_valid => p4_valid_1502, next_active_packet => next_active_packet_1553, next_pkt_with_priority => next_pkt_with_priority_1553); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_4_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity prioritySelect_Volatile is -- 
  port ( -- 
    down_counter : in  std_logic_vector(15 downto 0);
    active_packet : in  std_logic_vector(2 downto 0);
    pkt_with_priority : in  std_logic_vector(2 downto 0);
    p1_valid : in  std_logic_vector(0 downto 0);
    p2_valid : in  std_logic_vector(0 downto 0);
    p3_valid : in  std_logic_vector(0 downto 0);
    p4_valid : in  std_logic_vector(0 downto 0);
    next_active_packet : out  std_logic_vector(2 downto 0);
    next_pkt_with_priority : out  std_logic_vector(2 downto 0)-- 
  );
  -- 
end entity prioritySelect_Volatile;
architecture prioritySelect_Volatile_arch of prioritySelect_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(26-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal down_counter_buffer :  std_logic_vector(15 downto 0);
  signal active_packet_buffer :  std_logic_vector(2 downto 0);
  signal pkt_with_priority_buffer :  std_logic_vector(2 downto 0);
  signal p1_valid_buffer :  std_logic_vector(0 downto 0);
  signal p2_valid_buffer :  std_logic_vector(0 downto 0);
  signal p3_valid_buffer :  std_logic_vector(0 downto 0);
  signal p4_valid_buffer :  std_logic_vector(0 downto 0);
  -- output port buffer signals
  signal next_active_packet_buffer :  std_logic_vector(2 downto 0);
  signal next_pkt_with_priority_buffer :  std_logic_vector(2 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  down_counter_buffer <= down_counter;
  active_packet_buffer <= active_packet;
  pkt_with_priority_buffer <= pkt_with_priority;
  p1_valid_buffer <= p1_valid;
  p2_valid_buffer <= p2_valid;
  p3_valid_buffer <= p3_valid;
  p4_valid_buffer <= p4_valid;
  -- output handling  -------------------------------------------------------
  next_active_packet <= next_active_packet_buffer;
  next_pkt_with_priority <= next_pkt_with_priority_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_502_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_501_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_509_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_513_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_517_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_527_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_531_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_535_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_545_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_549_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_553_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_563_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_567_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_571_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_581_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_585_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_589_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_599_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_603_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_607_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_641_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_645_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_649_wire : std_logic_vector(0 downto 0);
    signal MUX_520_wire : std_logic_vector(0 downto 0);
    signal MUX_521_wire : std_logic_vector(0 downto 0);
    signal MUX_538_wire : std_logic_vector(0 downto 0);
    signal MUX_539_wire : std_logic_vector(0 downto 0);
    signal MUX_556_wire : std_logic_vector(2 downto 0);
    signal MUX_557_wire : std_logic_vector(2 downto 0);
    signal MUX_574_wire : std_logic_vector(0 downto 0);
    signal MUX_575_wire : std_logic_vector(0 downto 0);
    signal MUX_592_wire : std_logic_vector(2 downto 0);
    signal MUX_593_wire : std_logic_vector(2 downto 0);
    signal MUX_610_wire : std_logic_vector(0 downto 0);
    signal MUX_611_wire : std_logic_vector(0 downto 0);
    signal MUX_626_wire : std_logic_vector(2 downto 0);
    signal MUX_627_wire : std_logic_vector(2 downto 0);
    signal MUX_628_wire : std_logic_vector(2 downto 0);
    signal MUX_629_wire : std_logic_vector(2 downto 0);
    signal MUX_652_wire : std_logic_vector(2 downto 0);
    signal MUX_653_wire : std_logic_vector(2 downto 0);
    signal active_packet_priority_valid_541 : std_logic_vector(0 downto 0);
    signal check_pkt_4_505 : std_logic_vector(0 downto 0);
    signal d0_496 : std_logic_vector(0 downto 0);
    signal konst_494_wire_constant : std_logic_vector(15 downto 0);
    signal konst_500_wire_constant : std_logic_vector(2 downto 0);
    signal konst_508_wire_constant : std_logic_vector(2 downto 0);
    signal konst_512_wire_constant : std_logic_vector(2 downto 0);
    signal konst_516_wire_constant : std_logic_vector(2 downto 0);
    signal konst_526_wire_constant : std_logic_vector(2 downto 0);
    signal konst_530_wire_constant : std_logic_vector(2 downto 0);
    signal konst_534_wire_constant : std_logic_vector(2 downto 0);
    signal konst_544_wire_constant : std_logic_vector(2 downto 0);
    signal konst_546_wire_constant : std_logic_vector(2 downto 0);
    signal konst_548_wire_constant : std_logic_vector(2 downto 0);
    signal konst_550_wire_constant : std_logic_vector(2 downto 0);
    signal konst_552_wire_constant : std_logic_vector(2 downto 0);
    signal konst_554_wire_constant : std_logic_vector(2 downto 0);
    signal konst_555_wire_constant : std_logic_vector(2 downto 0);
    signal konst_562_wire_constant : std_logic_vector(2 downto 0);
    signal konst_566_wire_constant : std_logic_vector(2 downto 0);
    signal konst_570_wire_constant : std_logic_vector(2 downto 0);
    signal konst_580_wire_constant : std_logic_vector(2 downto 0);
    signal konst_582_wire_constant : std_logic_vector(2 downto 0);
    signal konst_584_wire_constant : std_logic_vector(2 downto 0);
    signal konst_586_wire_constant : std_logic_vector(2 downto 0);
    signal konst_588_wire_constant : std_logic_vector(2 downto 0);
    signal konst_590_wire_constant : std_logic_vector(2 downto 0);
    signal konst_591_wire_constant : std_logic_vector(2 downto 0);
    signal konst_598_wire_constant : std_logic_vector(2 downto 0);
    signal konst_602_wire_constant : std_logic_vector(2 downto 0);
    signal konst_606_wire_constant : std_logic_vector(2 downto 0);
    signal konst_616_wire_constant : std_logic_vector(2 downto 0);
    signal konst_625_wire_constant : std_logic_vector(2 downto 0);
    signal konst_640_wire_constant : std_logic_vector(2 downto 0);
    signal konst_642_wire_constant : std_logic_vector(2 downto 0);
    signal konst_644_wire_constant : std_logic_vector(2 downto 0);
    signal konst_646_wire_constant : std_logic_vector(2 downto 0);
    signal konst_648_wire_constant : std_logic_vector(2 downto 0);
    signal konst_650_wire_constant : std_logic_vector(2 downto 0);
    signal konst_651_wire_constant : std_logic_vector(2 downto 0);
    signal last_pkt_with_priority_595 : std_logic_vector(2 downto 0);
    signal last_pkt_with_priority_valid_613 : std_logic_vector(0 downto 0);
    signal next_to_pkt_with_priority_559 : std_logic_vector(2 downto 0);
    signal next_to_pkt_with_priority_valid_577 : std_logic_vector(0 downto 0);
    signal pkt_with_priority_valid_523 : std_logic_vector(0 downto 0);
    signal selected_packet_631 : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    konst_494_wire_constant <= "0000000000000000";
    konst_500_wire_constant <= "000";
    konst_508_wire_constant <= "001";
    konst_512_wire_constant <= "010";
    konst_516_wire_constant <= "011";
    konst_526_wire_constant <= "001";
    konst_530_wire_constant <= "010";
    konst_534_wire_constant <= "011";
    konst_544_wire_constant <= "001";
    konst_546_wire_constant <= "010";
    konst_548_wire_constant <= "010";
    konst_550_wire_constant <= "011";
    konst_552_wire_constant <= "011";
    konst_554_wire_constant <= "100";
    konst_555_wire_constant <= "001";
    konst_562_wire_constant <= "001";
    konst_566_wire_constant <= "010";
    konst_570_wire_constant <= "011";
    konst_580_wire_constant <= "001";
    konst_582_wire_constant <= "010";
    konst_584_wire_constant <= "010";
    konst_586_wire_constant <= "011";
    konst_588_wire_constant <= "011";
    konst_590_wire_constant <= "100";
    konst_591_wire_constant <= "001";
    konst_598_wire_constant <= "001";
    konst_602_wire_constant <= "010";
    konst_606_wire_constant <= "011";
    konst_616_wire_constant <= "100";
    konst_625_wire_constant <= "000";
    konst_640_wire_constant <= "001";
    konst_642_wire_constant <= "010";
    konst_644_wire_constant <= "010";
    konst_646_wire_constant <= "011";
    konst_648_wire_constant <= "011";
    konst_650_wire_constant <= "100";
    konst_651_wire_constant <= "001";
    -- flow-through select operator MUX_520_inst
    MUX_520_wire <= p3_valid_buffer when (EQ_u3_u1_517_wire(0) /=  '0') else p4_valid_buffer;
    -- flow-through select operator MUX_521_inst
    MUX_521_wire <= p2_valid_buffer when (EQ_u3_u1_513_wire(0) /=  '0') else MUX_520_wire;
    -- flow-through select operator MUX_522_inst
    pkt_with_priority_valid_523 <= p1_valid_buffer when (EQ_u3_u1_509_wire(0) /=  '0') else MUX_521_wire;
    -- flow-through select operator MUX_538_inst
    MUX_538_wire <= p3_valid_buffer when (EQ_u3_u1_535_wire(0) /=  '0') else p4_valid_buffer;
    -- flow-through select operator MUX_539_inst
    MUX_539_wire <= p2_valid_buffer when (EQ_u3_u1_531_wire(0) /=  '0') else MUX_538_wire;
    -- flow-through select operator MUX_540_inst
    active_packet_priority_valid_541 <= p1_valid_buffer when (EQ_u3_u1_527_wire(0) /=  '0') else MUX_539_wire;
    -- flow-through select operator MUX_556_inst
    MUX_556_wire <= konst_554_wire_constant when (EQ_u3_u1_553_wire(0) /=  '0') else konst_555_wire_constant;
    -- flow-through select operator MUX_557_inst
    MUX_557_wire <= konst_550_wire_constant when (EQ_u3_u1_549_wire(0) /=  '0') else MUX_556_wire;
    -- flow-through select operator MUX_558_inst
    next_to_pkt_with_priority_559 <= konst_546_wire_constant when (EQ_u3_u1_545_wire(0) /=  '0') else MUX_557_wire;
    -- flow-through select operator MUX_574_inst
    MUX_574_wire <= p3_valid_buffer when (EQ_u3_u1_571_wire(0) /=  '0') else p4_valid_buffer;
    -- flow-through select operator MUX_575_inst
    MUX_575_wire <= p2_valid_buffer when (EQ_u3_u1_567_wire(0) /=  '0') else MUX_574_wire;
    -- flow-through select operator MUX_576_inst
    next_to_pkt_with_priority_valid_577 <= p1_valid_buffer when (EQ_u3_u1_563_wire(0) /=  '0') else MUX_575_wire;
    -- flow-through select operator MUX_592_inst
    MUX_592_wire <= konst_590_wire_constant when (EQ_u3_u1_589_wire(0) /=  '0') else konst_591_wire_constant;
    -- flow-through select operator MUX_593_inst
    MUX_593_wire <= konst_586_wire_constant when (EQ_u3_u1_585_wire(0) /=  '0') else MUX_592_wire;
    -- flow-through select operator MUX_594_inst
    last_pkt_with_priority_595 <= konst_582_wire_constant when (EQ_u3_u1_581_wire(0) /=  '0') else MUX_593_wire;
    -- flow-through select operator MUX_610_inst
    MUX_610_wire <= p3_valid_buffer when (EQ_u3_u1_607_wire(0) /=  '0') else p4_valid_buffer;
    -- flow-through select operator MUX_611_inst
    MUX_611_wire <= p2_valid_buffer when (EQ_u3_u1_603_wire(0) /=  '0') else MUX_610_wire;
    -- flow-through select operator MUX_612_inst
    last_pkt_with_priority_valid_613 <= p1_valid_buffer when (EQ_u3_u1_599_wire(0) /=  '0') else MUX_611_wire;
    -- flow-through select operator MUX_626_inst
    MUX_626_wire <= active_packet_buffer when (active_packet_priority_valid_541(0) /=  '0') else konst_625_wire_constant;
    -- flow-through select operator MUX_627_inst
    MUX_627_wire <= last_pkt_with_priority_595 when (last_pkt_with_priority_valid_613(0) /=  '0') else MUX_626_wire;
    -- flow-through select operator MUX_628_inst
    MUX_628_wire <= next_to_pkt_with_priority_559 when (next_to_pkt_with_priority_valid_577(0) /=  '0') else MUX_627_wire;
    -- flow-through select operator MUX_629_inst
    MUX_629_wire <= pkt_with_priority_buffer when (pkt_with_priority_valid_523(0) /=  '0') else MUX_628_wire;
    -- flow-through select operator MUX_630_inst
    selected_packet_631 <= konst_616_wire_constant when (check_pkt_4_505(0) /=  '0') else MUX_629_wire;
    -- flow-through select operator MUX_636_inst
    next_active_packet_buffer <= selected_packet_631 when (d0_496(0) /=  '0') else active_packet_buffer;
    -- flow-through select operator MUX_652_inst
    MUX_652_wire <= konst_650_wire_constant when (EQ_u3_u1_649_wire(0) /=  '0') else konst_651_wire_constant;
    -- flow-through select operator MUX_653_inst
    MUX_653_wire <= konst_646_wire_constant when (EQ_u3_u1_645_wire(0) /=  '0') else MUX_652_wire;
    -- flow-through select operator MUX_654_inst
    next_pkt_with_priority_buffer <= konst_642_wire_constant when (EQ_u3_u1_641_wire(0) /=  '0') else MUX_653_wire;
    -- binary operator AND_u1_u1_502_inst
    process(d0_496, EQ_u3_u1_501_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_496, EQ_u3_u1_501_wire, tmp_var);
      AND_u1_u1_502_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_504_inst
    process(AND_u1_u1_502_wire, p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_502_wire, p4_valid_buffer, tmp_var);
      check_pkt_4_505 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_495_inst
    process(down_counter_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_buffer, konst_494_wire_constant, tmp_var);
      d0_496 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_501_inst
    process(active_packet_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_buffer, konst_500_wire_constant, tmp_var);
      EQ_u3_u1_501_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_509_inst
    process(pkt_with_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_with_priority_buffer, konst_508_wire_constant, tmp_var);
      EQ_u3_u1_509_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_513_inst
    process(pkt_with_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_with_priority_buffer, konst_512_wire_constant, tmp_var);
      EQ_u3_u1_513_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_517_inst
    process(pkt_with_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_with_priority_buffer, konst_516_wire_constant, tmp_var);
      EQ_u3_u1_517_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_527_inst
    process(active_packet_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_buffer, konst_526_wire_constant, tmp_var);
      EQ_u3_u1_527_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_531_inst
    process(active_packet_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_buffer, konst_530_wire_constant, tmp_var);
      EQ_u3_u1_531_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_535_inst
    process(active_packet_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_buffer, konst_534_wire_constant, tmp_var);
      EQ_u3_u1_535_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_545_inst
    process(pkt_with_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_with_priority_buffer, konst_544_wire_constant, tmp_var);
      EQ_u3_u1_545_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_549_inst
    process(pkt_with_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_with_priority_buffer, konst_548_wire_constant, tmp_var);
      EQ_u3_u1_549_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_553_inst
    process(pkt_with_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_with_priority_buffer, konst_552_wire_constant, tmp_var);
      EQ_u3_u1_553_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_563_inst
    process(next_to_pkt_with_priority_559) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_to_pkt_with_priority_559, konst_562_wire_constant, tmp_var);
      EQ_u3_u1_563_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_567_inst
    process(next_to_pkt_with_priority_559) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_to_pkt_with_priority_559, konst_566_wire_constant, tmp_var);
      EQ_u3_u1_567_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_571_inst
    process(next_to_pkt_with_priority_559) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_to_pkt_with_priority_559, konst_570_wire_constant, tmp_var);
      EQ_u3_u1_571_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_581_inst
    process(next_to_pkt_with_priority_559) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_to_pkt_with_priority_559, konst_580_wire_constant, tmp_var);
      EQ_u3_u1_581_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_585_inst
    process(next_to_pkt_with_priority_559) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_to_pkt_with_priority_559, konst_584_wire_constant, tmp_var);
      EQ_u3_u1_585_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_589_inst
    process(next_to_pkt_with_priority_559) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_to_pkt_with_priority_559, konst_588_wire_constant, tmp_var);
      EQ_u3_u1_589_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_599_inst
    process(last_pkt_with_priority_595) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last_pkt_with_priority_595, konst_598_wire_constant, tmp_var);
      EQ_u3_u1_599_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_603_inst
    process(last_pkt_with_priority_595) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last_pkt_with_priority_595, konst_602_wire_constant, tmp_var);
      EQ_u3_u1_603_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_607_inst
    process(last_pkt_with_priority_595) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last_pkt_with_priority_595, konst_606_wire_constant, tmp_var);
      EQ_u3_u1_607_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_641_inst
    process(next_active_packet_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_buffer, konst_640_wire_constant, tmp_var);
      EQ_u3_u1_641_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_645_inst
    process(next_active_packet_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_buffer, konst_644_wire_constant, tmp_var);
      EQ_u3_u1_645_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_649_inst
    process(next_active_packet_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_buffer, konst_648_wire_constant, tmp_var);
      EQ_u3_u1_649_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end prioritySelect_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_1_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_1_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_1_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_2_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_2_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_2_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_3_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_3_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_3_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_4_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_4_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_4_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_1_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_1_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_1_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_2_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_2_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_2_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_3_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_3_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_3_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_4_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_4_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_4_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- declarations related to module inputPort_1_Daemon
  component inputPort_1_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_1_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_1_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_1_Daemon
  signal inputPort_1_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_1_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_1_Daemon_start_req : std_logic;
  signal inputPort_1_Daemon_start_ack : std_logic;
  signal inputPort_1_Daemon_fin_req   : std_logic;
  signal inputPort_1_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_2_Daemon
  component inputPort_2_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_2_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_2_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_2_Daemon
  signal inputPort_2_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_2_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_2_Daemon_start_req : std_logic;
  signal inputPort_2_Daemon_start_ack : std_logic;
  signal inputPort_2_Daemon_fin_req   : std_logic;
  signal inputPort_2_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_3_Daemon
  component inputPort_3_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_3_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_3_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_3_Daemon
  signal inputPort_3_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_3_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_3_Daemon_start_req : std_logic;
  signal inputPort_3_Daemon_start_ack : std_logic;
  signal inputPort_3_Daemon_fin_req   : std_logic;
  signal inputPort_3_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_4_Daemon
  component inputPort_4_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_4_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_4_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_4_Daemon
  signal inputPort_4_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_4_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_4_Daemon_start_req : std_logic;
  signal inputPort_4_Daemon_start_ack : std_logic;
  signal inputPort_4_Daemon_fin_req   : std_logic;
  signal inputPort_4_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_1_Daemon
  component outputPort_1_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_1_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_1_Daemon
  signal outputPort_1_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_1_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_1_Daemon_start_req : std_logic;
  signal outputPort_1_Daemon_start_ack : std_logic;
  signal outputPort_1_Daemon_fin_req   : std_logic;
  signal outputPort_1_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_2_Daemon
  component outputPort_2_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_2_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_2_Daemon
  signal outputPort_2_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_2_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_2_Daemon_start_req : std_logic;
  signal outputPort_2_Daemon_start_ack : std_logic;
  signal outputPort_2_Daemon_fin_req   : std_logic;
  signal outputPort_2_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_3_Daemon
  component outputPort_3_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_3_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_3_Daemon
  signal outputPort_3_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_3_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_3_Daemon_start_req : std_logic;
  signal outputPort_3_Daemon_start_ack : std_logic;
  signal outputPort_3_Daemon_fin_req   : std_logic;
  signal outputPort_3_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_4_Daemon
  component outputPort_4_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_4_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_4_Daemon
  signal outputPort_4_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_4_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_4_Daemon_start_req : std_logic;
  signal outputPort_4_Daemon_start_ack : std_logic;
  signal outputPort_4_Daemon_fin_req   : std_logic;
  signal outputPort_4_Daemon_fin_ack : std_logic;
  -- declarations related to module prioritySelect
  -- aggregate signals for read from pipe in_data_1
  signal in_data_1_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_2
  signal in_data_2_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_3
  signal in_data_3_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_4
  signal in_data_4_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_1
  signal noblock_obuf_1_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_1
  signal noblock_obuf_1_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_2
  signal noblock_obuf_1_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_2
  signal noblock_obuf_1_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_3
  signal noblock_obuf_1_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_3
  signal noblock_obuf_1_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_4
  signal noblock_obuf_1_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_4
  signal noblock_obuf_1_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_1
  signal noblock_obuf_2_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_1
  signal noblock_obuf_2_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_2
  signal noblock_obuf_2_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_2
  signal noblock_obuf_2_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_3
  signal noblock_obuf_2_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_3
  signal noblock_obuf_2_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_4
  signal noblock_obuf_2_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_4
  signal noblock_obuf_2_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_1
  signal noblock_obuf_3_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_1
  signal noblock_obuf_3_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_2
  signal noblock_obuf_3_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_2
  signal noblock_obuf_3_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_3
  signal noblock_obuf_3_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_3
  signal noblock_obuf_3_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_4
  signal noblock_obuf_3_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_4
  signal noblock_obuf_3_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_1
  signal noblock_obuf_4_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_1
  signal noblock_obuf_4_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_2
  signal noblock_obuf_4_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_2
  signal noblock_obuf_4_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_3
  signal noblock_obuf_4_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_3
  signal noblock_obuf_4_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_4
  signal noblock_obuf_4_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_4
  signal noblock_obuf_4_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_1
  signal out_data_1_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_2
  signal out_data_2_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_3
  signal out_data_3_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_4
  signal out_data_4_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module inputPort_1_Daemon
  inputPort_1_Daemon_instance:inputPort_1_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_1_Daemon_start_req,
      start_ack => inputPort_1_Daemon_start_ack,
      fin_req => inputPort_1_Daemon_fin_req,
      fin_ack => inputPort_1_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_1_pipe_read_req => in_data_1_pipe_read_req(0 downto 0),
      in_data_1_pipe_read_ack => in_data_1_pipe_read_ack(0 downto 0),
      in_data_1_pipe_read_data => in_data_1_pipe_read_data(31 downto 0),
      noblock_obuf_1_1_pipe_write_req => noblock_obuf_1_1_pipe_write_req(0 downto 0),
      noblock_obuf_1_1_pipe_write_ack => noblock_obuf_1_1_pipe_write_ack(0 downto 0),
      noblock_obuf_1_1_pipe_write_data => noblock_obuf_1_1_pipe_write_data(32 downto 0),
      noblock_obuf_1_3_pipe_write_req => noblock_obuf_1_3_pipe_write_req(0 downto 0),
      noblock_obuf_1_3_pipe_write_ack => noblock_obuf_1_3_pipe_write_ack(0 downto 0),
      noblock_obuf_1_3_pipe_write_data => noblock_obuf_1_3_pipe_write_data(32 downto 0),
      noblock_obuf_1_4_pipe_write_req => noblock_obuf_1_4_pipe_write_req(0 downto 0),
      noblock_obuf_1_4_pipe_write_ack => noblock_obuf_1_4_pipe_write_ack(0 downto 0),
      noblock_obuf_1_4_pipe_write_data => noblock_obuf_1_4_pipe_write_data(32 downto 0),
      noblock_obuf_1_2_pipe_write_req => noblock_obuf_1_2_pipe_write_req(0 downto 0),
      noblock_obuf_1_2_pipe_write_ack => noblock_obuf_1_2_pipe_write_ack(0 downto 0),
      noblock_obuf_1_2_pipe_write_data => noblock_obuf_1_2_pipe_write_data(32 downto 0),
      tag_in => inputPort_1_Daemon_tag_in,
      tag_out => inputPort_1_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_1_Daemon_tag_in <= (others => '0');
  inputPort_1_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_1_Daemon_start_req, start_ack => inputPort_1_Daemon_start_ack,  fin_req => inputPort_1_Daemon_fin_req,  fin_ack => inputPort_1_Daemon_fin_ack);
  -- module inputPort_2_Daemon
  inputPort_2_Daemon_instance:inputPort_2_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_2_Daemon_start_req,
      start_ack => inputPort_2_Daemon_start_ack,
      fin_req => inputPort_2_Daemon_fin_req,
      fin_ack => inputPort_2_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_2_pipe_read_req => in_data_2_pipe_read_req(0 downto 0),
      in_data_2_pipe_read_ack => in_data_2_pipe_read_ack(0 downto 0),
      in_data_2_pipe_read_data => in_data_2_pipe_read_data(31 downto 0),
      noblock_obuf_2_1_pipe_write_req => noblock_obuf_2_1_pipe_write_req(0 downto 0),
      noblock_obuf_2_1_pipe_write_ack => noblock_obuf_2_1_pipe_write_ack(0 downto 0),
      noblock_obuf_2_1_pipe_write_data => noblock_obuf_2_1_pipe_write_data(32 downto 0),
      noblock_obuf_2_2_pipe_write_req => noblock_obuf_2_2_pipe_write_req(0 downto 0),
      noblock_obuf_2_2_pipe_write_ack => noblock_obuf_2_2_pipe_write_ack(0 downto 0),
      noblock_obuf_2_2_pipe_write_data => noblock_obuf_2_2_pipe_write_data(32 downto 0),
      noblock_obuf_2_3_pipe_write_req => noblock_obuf_2_3_pipe_write_req(0 downto 0),
      noblock_obuf_2_3_pipe_write_ack => noblock_obuf_2_3_pipe_write_ack(0 downto 0),
      noblock_obuf_2_3_pipe_write_data => noblock_obuf_2_3_pipe_write_data(32 downto 0),
      noblock_obuf_2_4_pipe_write_req => noblock_obuf_2_4_pipe_write_req(0 downto 0),
      noblock_obuf_2_4_pipe_write_ack => noblock_obuf_2_4_pipe_write_ack(0 downto 0),
      noblock_obuf_2_4_pipe_write_data => noblock_obuf_2_4_pipe_write_data(32 downto 0),
      tag_in => inputPort_2_Daemon_tag_in,
      tag_out => inputPort_2_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_2_Daemon_tag_in <= (others => '0');
  inputPort_2_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_2_Daemon_start_req, start_ack => inputPort_2_Daemon_start_ack,  fin_req => inputPort_2_Daemon_fin_req,  fin_ack => inputPort_2_Daemon_fin_ack);
  -- module inputPort_3_Daemon
  inputPort_3_Daemon_instance:inputPort_3_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_3_Daemon_start_req,
      start_ack => inputPort_3_Daemon_start_ack,
      fin_req => inputPort_3_Daemon_fin_req,
      fin_ack => inputPort_3_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_3_pipe_read_req => in_data_3_pipe_read_req(0 downto 0),
      in_data_3_pipe_read_ack => in_data_3_pipe_read_ack(0 downto 0),
      in_data_3_pipe_read_data => in_data_3_pipe_read_data(31 downto 0),
      noblock_obuf_3_2_pipe_write_req => noblock_obuf_3_2_pipe_write_req(0 downto 0),
      noblock_obuf_3_2_pipe_write_ack => noblock_obuf_3_2_pipe_write_ack(0 downto 0),
      noblock_obuf_3_2_pipe_write_data => noblock_obuf_3_2_pipe_write_data(32 downto 0),
      noblock_obuf_3_3_pipe_write_req => noblock_obuf_3_3_pipe_write_req(0 downto 0),
      noblock_obuf_3_3_pipe_write_ack => noblock_obuf_3_3_pipe_write_ack(0 downto 0),
      noblock_obuf_3_3_pipe_write_data => noblock_obuf_3_3_pipe_write_data(32 downto 0),
      noblock_obuf_3_4_pipe_write_req => noblock_obuf_3_4_pipe_write_req(0 downto 0),
      noblock_obuf_3_4_pipe_write_ack => noblock_obuf_3_4_pipe_write_ack(0 downto 0),
      noblock_obuf_3_4_pipe_write_data => noblock_obuf_3_4_pipe_write_data(32 downto 0),
      noblock_obuf_3_1_pipe_write_req => noblock_obuf_3_1_pipe_write_req(0 downto 0),
      noblock_obuf_3_1_pipe_write_ack => noblock_obuf_3_1_pipe_write_ack(0 downto 0),
      noblock_obuf_3_1_pipe_write_data => noblock_obuf_3_1_pipe_write_data(32 downto 0),
      tag_in => inputPort_3_Daemon_tag_in,
      tag_out => inputPort_3_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_3_Daemon_tag_in <= (others => '0');
  inputPort_3_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_3_Daemon_start_req, start_ack => inputPort_3_Daemon_start_ack,  fin_req => inputPort_3_Daemon_fin_req,  fin_ack => inputPort_3_Daemon_fin_ack);
  -- module inputPort_4_Daemon
  inputPort_4_Daemon_instance:inputPort_4_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_4_Daemon_start_req,
      start_ack => inputPort_4_Daemon_start_ack,
      fin_req => inputPort_4_Daemon_fin_req,
      fin_ack => inputPort_4_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_4_pipe_read_req => in_data_4_pipe_read_req(0 downto 0),
      in_data_4_pipe_read_ack => in_data_4_pipe_read_ack(0 downto 0),
      in_data_4_pipe_read_data => in_data_4_pipe_read_data(31 downto 0),
      noblock_obuf_4_1_pipe_write_req => noblock_obuf_4_1_pipe_write_req(0 downto 0),
      noblock_obuf_4_1_pipe_write_ack => noblock_obuf_4_1_pipe_write_ack(0 downto 0),
      noblock_obuf_4_1_pipe_write_data => noblock_obuf_4_1_pipe_write_data(32 downto 0),
      noblock_obuf_4_2_pipe_write_req => noblock_obuf_4_2_pipe_write_req(0 downto 0),
      noblock_obuf_4_2_pipe_write_ack => noblock_obuf_4_2_pipe_write_ack(0 downto 0),
      noblock_obuf_4_2_pipe_write_data => noblock_obuf_4_2_pipe_write_data(32 downto 0),
      noblock_obuf_4_3_pipe_write_req => noblock_obuf_4_3_pipe_write_req(0 downto 0),
      noblock_obuf_4_3_pipe_write_ack => noblock_obuf_4_3_pipe_write_ack(0 downto 0),
      noblock_obuf_4_3_pipe_write_data => noblock_obuf_4_3_pipe_write_data(32 downto 0),
      noblock_obuf_4_4_pipe_write_req => noblock_obuf_4_4_pipe_write_req(0 downto 0),
      noblock_obuf_4_4_pipe_write_ack => noblock_obuf_4_4_pipe_write_ack(0 downto 0),
      noblock_obuf_4_4_pipe_write_data => noblock_obuf_4_4_pipe_write_data(32 downto 0),
      tag_in => inputPort_4_Daemon_tag_in,
      tag_out => inputPort_4_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_4_Daemon_tag_in <= (others => '0');
  inputPort_4_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_4_Daemon_start_req, start_ack => inputPort_4_Daemon_start_ack,  fin_req => inputPort_4_Daemon_fin_req,  fin_ack => inputPort_4_Daemon_fin_ack);
  -- module outputPort_1_Daemon
  outputPort_1_Daemon_instance:outputPort_1_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_1_Daemon_start_req,
      start_ack => outputPort_1_Daemon_start_ack,
      fin_req => outputPort_1_Daemon_fin_req,
      fin_ack => outputPort_1_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_1_pipe_read_req => noblock_obuf_1_1_pipe_read_req(0 downto 0),
      noblock_obuf_1_1_pipe_read_ack => noblock_obuf_1_1_pipe_read_ack(0 downto 0),
      noblock_obuf_1_1_pipe_read_data => noblock_obuf_1_1_pipe_read_data(32 downto 0),
      noblock_obuf_2_1_pipe_read_req => noblock_obuf_2_1_pipe_read_req(0 downto 0),
      noblock_obuf_2_1_pipe_read_ack => noblock_obuf_2_1_pipe_read_ack(0 downto 0),
      noblock_obuf_2_1_pipe_read_data => noblock_obuf_2_1_pipe_read_data(32 downto 0),
      noblock_obuf_4_1_pipe_read_req => noblock_obuf_4_1_pipe_read_req(0 downto 0),
      noblock_obuf_4_1_pipe_read_ack => noblock_obuf_4_1_pipe_read_ack(0 downto 0),
      noblock_obuf_4_1_pipe_read_data => noblock_obuf_4_1_pipe_read_data(32 downto 0),
      noblock_obuf_3_1_pipe_read_req => noblock_obuf_3_1_pipe_read_req(0 downto 0),
      noblock_obuf_3_1_pipe_read_ack => noblock_obuf_3_1_pipe_read_ack(0 downto 0),
      noblock_obuf_3_1_pipe_read_data => noblock_obuf_3_1_pipe_read_data(32 downto 0),
      out_data_1_pipe_write_req => out_data_1_pipe_write_req(0 downto 0),
      out_data_1_pipe_write_ack => out_data_1_pipe_write_ack(0 downto 0),
      out_data_1_pipe_write_data => out_data_1_pipe_write_data(31 downto 0),
      tag_in => outputPort_1_Daemon_tag_in,
      tag_out => outputPort_1_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_1_Daemon_tag_in <= (others => '0');
  outputPort_1_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_1_Daemon_start_req, start_ack => outputPort_1_Daemon_start_ack,  fin_req => outputPort_1_Daemon_fin_req,  fin_ack => outputPort_1_Daemon_fin_ack);
  -- module outputPort_2_Daemon
  outputPort_2_Daemon_instance:outputPort_2_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_2_Daemon_start_req,
      start_ack => outputPort_2_Daemon_start_ack,
      fin_req => outputPort_2_Daemon_fin_req,
      fin_ack => outputPort_2_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_2_pipe_read_req => noblock_obuf_1_2_pipe_read_req(0 downto 0),
      noblock_obuf_1_2_pipe_read_ack => noblock_obuf_1_2_pipe_read_ack(0 downto 0),
      noblock_obuf_1_2_pipe_read_data => noblock_obuf_1_2_pipe_read_data(32 downto 0),
      noblock_obuf_3_2_pipe_read_req => noblock_obuf_3_2_pipe_read_req(0 downto 0),
      noblock_obuf_3_2_pipe_read_ack => noblock_obuf_3_2_pipe_read_ack(0 downto 0),
      noblock_obuf_3_2_pipe_read_data => noblock_obuf_3_2_pipe_read_data(32 downto 0),
      noblock_obuf_4_2_pipe_read_req => noblock_obuf_4_2_pipe_read_req(0 downto 0),
      noblock_obuf_4_2_pipe_read_ack => noblock_obuf_4_2_pipe_read_ack(0 downto 0),
      noblock_obuf_4_2_pipe_read_data => noblock_obuf_4_2_pipe_read_data(32 downto 0),
      noblock_obuf_2_2_pipe_read_req => noblock_obuf_2_2_pipe_read_req(0 downto 0),
      noblock_obuf_2_2_pipe_read_ack => noblock_obuf_2_2_pipe_read_ack(0 downto 0),
      noblock_obuf_2_2_pipe_read_data => noblock_obuf_2_2_pipe_read_data(32 downto 0),
      out_data_2_pipe_write_req => out_data_2_pipe_write_req(0 downto 0),
      out_data_2_pipe_write_ack => out_data_2_pipe_write_ack(0 downto 0),
      out_data_2_pipe_write_data => out_data_2_pipe_write_data(31 downto 0),
      tag_in => outputPort_2_Daemon_tag_in,
      tag_out => outputPort_2_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_2_Daemon_tag_in <= (others => '0');
  outputPort_2_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_2_Daemon_start_req, start_ack => outputPort_2_Daemon_start_ack,  fin_req => outputPort_2_Daemon_fin_req,  fin_ack => outputPort_2_Daemon_fin_ack);
  -- module outputPort_3_Daemon
  outputPort_3_Daemon_instance:outputPort_3_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_3_Daemon_start_req,
      start_ack => outputPort_3_Daemon_start_ack,
      fin_req => outputPort_3_Daemon_fin_req,
      fin_ack => outputPort_3_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_3_pipe_read_req => noblock_obuf_1_3_pipe_read_req(0 downto 0),
      noblock_obuf_1_3_pipe_read_ack => noblock_obuf_1_3_pipe_read_ack(0 downto 0),
      noblock_obuf_1_3_pipe_read_data => noblock_obuf_1_3_pipe_read_data(32 downto 0),
      noblock_obuf_3_3_pipe_read_req => noblock_obuf_3_3_pipe_read_req(0 downto 0),
      noblock_obuf_3_3_pipe_read_ack => noblock_obuf_3_3_pipe_read_ack(0 downto 0),
      noblock_obuf_3_3_pipe_read_data => noblock_obuf_3_3_pipe_read_data(32 downto 0),
      noblock_obuf_2_3_pipe_read_req => noblock_obuf_2_3_pipe_read_req(0 downto 0),
      noblock_obuf_2_3_pipe_read_ack => noblock_obuf_2_3_pipe_read_ack(0 downto 0),
      noblock_obuf_2_3_pipe_read_data => noblock_obuf_2_3_pipe_read_data(32 downto 0),
      noblock_obuf_4_3_pipe_read_req => noblock_obuf_4_3_pipe_read_req(0 downto 0),
      noblock_obuf_4_3_pipe_read_ack => noblock_obuf_4_3_pipe_read_ack(0 downto 0),
      noblock_obuf_4_3_pipe_read_data => noblock_obuf_4_3_pipe_read_data(32 downto 0),
      out_data_3_pipe_write_req => out_data_3_pipe_write_req(0 downto 0),
      out_data_3_pipe_write_ack => out_data_3_pipe_write_ack(0 downto 0),
      out_data_3_pipe_write_data => out_data_3_pipe_write_data(31 downto 0),
      tag_in => outputPort_3_Daemon_tag_in,
      tag_out => outputPort_3_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_3_Daemon_tag_in <= (others => '0');
  outputPort_3_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_3_Daemon_start_req, start_ack => outputPort_3_Daemon_start_ack,  fin_req => outputPort_3_Daemon_fin_req,  fin_ack => outputPort_3_Daemon_fin_ack);
  -- module outputPort_4_Daemon
  outputPort_4_Daemon_instance:outputPort_4_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_4_Daemon_start_req,
      start_ack => outputPort_4_Daemon_start_ack,
      fin_req => outputPort_4_Daemon_fin_req,
      fin_ack => outputPort_4_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_4_pipe_read_req => noblock_obuf_1_4_pipe_read_req(0 downto 0),
      noblock_obuf_1_4_pipe_read_ack => noblock_obuf_1_4_pipe_read_ack(0 downto 0),
      noblock_obuf_1_4_pipe_read_data => noblock_obuf_1_4_pipe_read_data(32 downto 0),
      noblock_obuf_3_4_pipe_read_req => noblock_obuf_3_4_pipe_read_req(0 downto 0),
      noblock_obuf_3_4_pipe_read_ack => noblock_obuf_3_4_pipe_read_ack(0 downto 0),
      noblock_obuf_3_4_pipe_read_data => noblock_obuf_3_4_pipe_read_data(32 downto 0),
      noblock_obuf_2_4_pipe_read_req => noblock_obuf_2_4_pipe_read_req(0 downto 0),
      noblock_obuf_2_4_pipe_read_ack => noblock_obuf_2_4_pipe_read_ack(0 downto 0),
      noblock_obuf_2_4_pipe_read_data => noblock_obuf_2_4_pipe_read_data(32 downto 0),
      noblock_obuf_4_4_pipe_read_req => noblock_obuf_4_4_pipe_read_req(0 downto 0),
      noblock_obuf_4_4_pipe_read_ack => noblock_obuf_4_4_pipe_read_ack(0 downto 0),
      noblock_obuf_4_4_pipe_read_data => noblock_obuf_4_4_pipe_read_data(32 downto 0),
      out_data_4_pipe_write_req => out_data_4_pipe_write_req(0 downto 0),
      out_data_4_pipe_write_ack => out_data_4_pipe_write_ack(0 downto 0),
      out_data_4_pipe_write_data => out_data_4_pipe_write_data(31 downto 0),
      tag_in => outputPort_4_Daemon_tag_in,
      tag_out => outputPort_4_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_4_Daemon_tag_in <= (others => '0');
  outputPort_4_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_4_Daemon_start_req, start_ack => outputPort_4_Daemon_start_ack,  fin_req => outputPort_4_Daemon_fin_req,  fin_ack => outputPort_4_Daemon_fin_ack);
  in_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_1_pipe_read_req,
      read_ack => in_data_1_pipe_read_ack,
      read_data => in_data_1_pipe_read_data,
      write_req => in_data_1_pipe_write_req,
      write_ack => in_data_1_pipe_write_ack,
      write_data => in_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_2_pipe_read_req,
      read_ack => in_data_2_pipe_read_ack,
      read_data => in_data_2_pipe_read_data,
      write_req => in_data_2_pipe_write_req,
      write_ack => in_data_2_pipe_write_ack,
      write_data => in_data_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_3_pipe_read_req,
      read_ack => in_data_3_pipe_read_ack,
      read_data => in_data_3_pipe_read_data,
      write_req => in_data_3_pipe_write_req,
      write_ack => in_data_3_pipe_write_ack,
      write_data => in_data_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_4_pipe_read_req,
      read_ack => in_data_4_pipe_read_ack,
      read_data => in_data_4_pipe_read_data,
      write_req => in_data_4_pipe_write_req,
      write_ack => in_data_4_pipe_write_ack,
      write_data => in_data_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_1_pipe_read_req,
      read_ack => noblock_obuf_1_1_pipe_read_ack,
      read_data => noblock_obuf_1_1_pipe_read_data,
      write_req => noblock_obuf_1_1_pipe_write_req,
      write_ack => noblock_obuf_1_1_pipe_write_ack,
      write_data => noblock_obuf_1_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_2_pipe_read_req,
      read_ack => noblock_obuf_1_2_pipe_read_ack,
      read_data => noblock_obuf_1_2_pipe_read_data,
      write_req => noblock_obuf_1_2_pipe_write_req,
      write_ack => noblock_obuf_1_2_pipe_write_ack,
      write_data => noblock_obuf_1_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_3_pipe_read_req,
      read_ack => noblock_obuf_1_3_pipe_read_ack,
      read_data => noblock_obuf_1_3_pipe_read_data,
      write_req => noblock_obuf_1_3_pipe_write_req,
      write_ack => noblock_obuf_1_3_pipe_write_ack,
      write_data => noblock_obuf_1_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_4_pipe_read_req,
      read_ack => noblock_obuf_1_4_pipe_read_ack,
      read_data => noblock_obuf_1_4_pipe_read_data,
      write_req => noblock_obuf_1_4_pipe_write_req,
      write_ack => noblock_obuf_1_4_pipe_write_ack,
      write_data => noblock_obuf_1_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_1_pipe_read_req,
      read_ack => noblock_obuf_2_1_pipe_read_ack,
      read_data => noblock_obuf_2_1_pipe_read_data,
      write_req => noblock_obuf_2_1_pipe_write_req,
      write_ack => noblock_obuf_2_1_pipe_write_ack,
      write_data => noblock_obuf_2_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_2_pipe_read_req,
      read_ack => noblock_obuf_2_2_pipe_read_ack,
      read_data => noblock_obuf_2_2_pipe_read_data,
      write_req => noblock_obuf_2_2_pipe_write_req,
      write_ack => noblock_obuf_2_2_pipe_write_ack,
      write_data => noblock_obuf_2_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_3_pipe_read_req,
      read_ack => noblock_obuf_2_3_pipe_read_ack,
      read_data => noblock_obuf_2_3_pipe_read_data,
      write_req => noblock_obuf_2_3_pipe_write_req,
      write_ack => noblock_obuf_2_3_pipe_write_ack,
      write_data => noblock_obuf_2_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_4_pipe_read_req,
      read_ack => noblock_obuf_2_4_pipe_read_ack,
      read_data => noblock_obuf_2_4_pipe_read_data,
      write_req => noblock_obuf_2_4_pipe_write_req,
      write_ack => noblock_obuf_2_4_pipe_write_ack,
      write_data => noblock_obuf_2_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_1_pipe_read_req,
      read_ack => noblock_obuf_3_1_pipe_read_ack,
      read_data => noblock_obuf_3_1_pipe_read_data,
      write_req => noblock_obuf_3_1_pipe_write_req,
      write_ack => noblock_obuf_3_1_pipe_write_ack,
      write_data => noblock_obuf_3_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_2_pipe_read_req,
      read_ack => noblock_obuf_3_2_pipe_read_ack,
      read_data => noblock_obuf_3_2_pipe_read_data,
      write_req => noblock_obuf_3_2_pipe_write_req,
      write_ack => noblock_obuf_3_2_pipe_write_ack,
      write_data => noblock_obuf_3_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_3_pipe_read_req,
      read_ack => noblock_obuf_3_3_pipe_read_ack,
      read_data => noblock_obuf_3_3_pipe_read_data,
      write_req => noblock_obuf_3_3_pipe_write_req,
      write_ack => noblock_obuf_3_3_pipe_write_ack,
      write_data => noblock_obuf_3_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_4_pipe_read_req,
      read_ack => noblock_obuf_3_4_pipe_read_ack,
      read_data => noblock_obuf_3_4_pipe_read_data,
      write_req => noblock_obuf_3_4_pipe_write_req,
      write_ack => noblock_obuf_3_4_pipe_write_ack,
      write_data => noblock_obuf_3_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_1_pipe_read_req,
      read_ack => noblock_obuf_4_1_pipe_read_ack,
      read_data => noblock_obuf_4_1_pipe_read_data,
      write_req => noblock_obuf_4_1_pipe_write_req,
      write_ack => noblock_obuf_4_1_pipe_write_ack,
      write_data => noblock_obuf_4_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_2_pipe_read_req,
      read_ack => noblock_obuf_4_2_pipe_read_ack,
      read_data => noblock_obuf_4_2_pipe_read_data,
      write_req => noblock_obuf_4_2_pipe_write_req,
      write_ack => noblock_obuf_4_2_pipe_write_ack,
      write_data => noblock_obuf_4_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_3_pipe_read_req,
      read_ack => noblock_obuf_4_3_pipe_read_ack,
      read_data => noblock_obuf_4_3_pipe_read_data,
      write_req => noblock_obuf_4_3_pipe_write_req,
      write_ack => noblock_obuf_4_3_pipe_write_ack,
      write_data => noblock_obuf_4_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_4_pipe_read_req,
      read_ack => noblock_obuf_4_4_pipe_read_ack,
      read_data => noblock_obuf_4_4_pipe_read_data,
      write_req => noblock_obuf_4_4_pipe_write_req,
      write_ack => noblock_obuf_4_4_pipe_write_ack,
      write_data => noblock_obuf_4_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_1_pipe_read_req,
      read_ack => out_data_1_pipe_read_ack,
      read_data => out_data_1_pipe_read_data,
      write_req => out_data_1_pipe_write_req,
      write_ack => out_data_1_pipe_write_ack,
      write_data => out_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_2_pipe_read_req,
      read_ack => out_data_2_pipe_read_ack,
      read_data => out_data_2_pipe_read_data,
      write_req => out_data_2_pipe_write_req,
      write_ack => out_data_2_pipe_write_ack,
      write_data => out_data_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_3_pipe_read_req,
      read_ack => out_data_3_pipe_read_ack,
      read_data => out_data_3_pipe_read_data,
      write_req => out_data_3_pipe_write_req,
      write_ack => out_data_3_pipe_write_ack,
      write_data => out_data_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_4_pipe_read_req,
      read_ack => out_data_4_pipe_read_ack,
      read_data => out_data_4_pipe_read_data,
      write_req => out_data_4_pipe_write_req,
      write_ack => out_data_4_pipe_write_ack,
      write_data => out_data_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- 
end ahir_system_arch;
